
//------> /hd/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /hd/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   saranyuc@rsg24.stanford.edu
//  Generated date: Wed Apr  8 16:36:33 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    aqed_top_core
// ------------------------------------------------------------------


module aqed_top_core (
  clk, clk_en, reset, bmc_in_rsc_dat, bmc_v_rsc_dat, original_rsc_dat, duplicate_rsc_dat,
      acc_out_rsc_dat, acc_out_v_rsc_dat, acc_out_rdy_rsc_dat, return_aqed_out_rsc_dat,
      return_aqed_out_v_rsc_dat, return_qed_done_rsc_dat, return_qed_check_rsc_dat,
      return_orig_issued_rsc_dat, return_orig_done_rsc_dat
);
  input clk;
  input clk_en;
  input reset;
  input [15:0] bmc_in_rsc_dat;
  input bmc_v_rsc_dat;
  input original_rsc_dat;
  input duplicate_rsc_dat;
  input [15:0] acc_out_rsc_dat;
  input acc_out_v_rsc_dat;
  input acc_out_rdy_rsc_dat;
  output [15:0] return_aqed_out_rsc_dat;
  output return_aqed_out_v_rsc_dat;
  output return_qed_done_rsc_dat;
  output return_qed_check_rsc_dat;
  output return_orig_issued_rsc_dat;
  output return_orig_done_rsc_dat;


  // Interconnect Declarations
  wire [15:0] bmc_in_rsci_idat;
  wire bmc_v_rsci_idat;
  wire original_rsci_idat;
  wire duplicate_rsci_idat;
  wire [15:0] acc_out_rsci_idat;
  wire acc_out_v_rsci_idat;
  wire acc_out_rdy_rsci_idat;
  reg [15:0] return_aqed_out_rsci_idat;
  reg return_aqed_out_v_rsci_idat;
  wire aqed_out_if_aif_4_equal_tmp;
  wire aqed_out_if_aif_1_equal_tmp;
  wire aqed_out_if_aqed_out_if_and_1_tmp;
  wire aqed_in_if_issue_dup_aif_1_aif_equal_tmp;
  wire state_dup_issued_sva_mx0;
  wire state_orig_issued_sva_dfm_1_mx0;
  wire aqed_in_if_issue_orig_land_lpi_1_dfm_1;
  reg state_orig_issued_sva;
  reg state_dup_issued_sva;
  reg state_qed_done_sva;
  reg reg_state_orig_done_cse;
  reg reg_state_qed_check_cse;
  wire and_9_cse;
  wire or_15_cse;
  wire mux_3_cse;
  wire state_out_count_and_cse;
  wire mux_1_itm;
  reg [15:0] state_orig_sva;
  reg [15:0] state_orig_in_sva;
  reg [15:0] state_orig_out_sva;
  reg [15:0] state_dup_in_sva;
  reg [15:0] state_in_count_sva;
  wire [16:0] nl_state_in_count_sva;
  reg [15:0] state_out_count_sva;
  wire [16:0] nl_state_out_count_sva;
  wire [15:0] state_orig_in_sva_dfm_1_mx0;
  wire [15:0] state_dup_in_sva_dfm_1_mx1;
  wire and_dcpl_10;
  wire mux_5_cse;
  wire aqed_out_if_if_2_acc_itm_16_1;

  wire[15:0] aqed_out_if_mux_2_nl;
  wire[0:0] aqed_out_if_if_aqed_out_if_if_and_1_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] nor_4_nl;
  wire[16:0] aqed_out_if_aelse_acc_nl;
  wire[18:0] nl_aqed_out_if_aelse_acc_nl;
  wire[0:0] and_6_nl;
  wire[15:0] state_in_count_mux_1_nl;
  wire[0:0] nand_3_nl;
  wire[16:0] aqed_out_if_if_2_acc_nl;
  wire[18:0] nl_aqed_out_if_if_2_acc_nl;
  wire[0:0] aqed_in_if_aqed_in_if_or_2_nl;
  wire[0:0] aqed_in_if_aqed_in_if_or_3_nl;
  wire[0:0] and_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_return_qed_done_rsci_idat;
  assign nl_return_qed_done_rsci_idat = state_qed_done_sva;
  wire [0:0] nl_return_qed_check_rsci_idat;
  assign nl_return_qed_check_rsci_idat = reg_state_qed_check_cse;
  wire [0:0] nl_return_orig_issued_rsci_idat;
  assign nl_return_orig_issued_rsci_idat = state_orig_issued_sva;
  wire [0:0] nl_return_orig_done_rsci_idat;
  assign nl_return_orig_done_rsci_idat = reg_state_orig_done_cse;
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd16)) bmc_in_rsci (
      .dat(bmc_in_rsc_dat),
      .idat(bmc_in_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd1)) bmc_v_rsci (
      .dat(bmc_v_rsc_dat),
      .idat(bmc_v_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd1)) original_rsci (
      .dat(original_rsc_dat),
      .idat(original_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd1)) duplicate_rsci (
      .dat(duplicate_rsc_dat),
      .idat(duplicate_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd16)) acc_out_rsci (
      .dat(acc_out_rsc_dat),
      .idat(acc_out_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd1)) acc_out_v_rsci (
      .dat(acc_out_v_rsc_dat),
      .idat(acc_out_v_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd1)) acc_out_rdy_rsci (
      .dat(acc_out_rdy_rsc_dat),
      .idat(acc_out_rdy_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd8),
  .width(32'sd16)) return_aqed_out_rsci (
      .idat(return_aqed_out_rsci_idat),
      .dat(return_aqed_out_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd9),
  .width(32'sd1)) return_aqed_out_v_rsci (
      .idat(return_aqed_out_v_rsci_idat),
      .dat(return_aqed_out_v_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd10),
  .width(32'sd1)) return_qed_done_rsci (
      .idat(nl_return_qed_done_rsci_idat[0:0]),
      .dat(return_qed_done_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd11),
  .width(32'sd1)) return_qed_check_rsci (
      .idat(nl_return_qed_check_rsci_idat[0:0]),
      .dat(return_qed_check_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd12),
  .width(32'sd1)) return_orig_issued_rsci (
      .idat(nl_return_orig_issued_rsci_idat[0:0]),
      .dat(return_orig_issued_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd13),
  .width(32'sd1)) return_orig_done_rsci (
      .idat(nl_return_orig_done_rsci_idat[0:0]),
      .dat(return_orig_done_rsc_dat)
    );
  assign and_9_cse = bmc_v_rsci_idat & original_rsci_idat;
  assign or_15_cse = and_9_cse | state_orig_issued_sva;
  assign state_out_count_and_cse = clk_en & aqed_out_if_aqed_out_if_and_1_tmp;
  assign aqed_out_if_aif_1_equal_tmp = state_out_count_sva == state_orig_in_sva_dfm_1_mx0;
  assign state_orig_in_sva_dfm_1_mx0 = MUX_v_16_2_2(state_in_count_sva, state_orig_in_sva,
      state_orig_issued_sva);
  assign and_6_nl = aqed_in_if_issue_dup_aif_1_aif_equal_tmp & bmc_v_rsci_idat;
  assign mux_3_cse = MUX_s_1_2_2(and_9_cse, (and_6_nl), state_orig_issued_sva);
  assign state_in_count_mux_1_nl = MUX_v_16_2_2(state_in_count_sva, state_dup_in_sva,
      state_dup_issued_sva);
  assign aqed_out_if_aif_4_equal_tmp = state_out_count_sva == (state_in_count_mux_1_nl);
  assign mux_5_cse = MUX_s_1_2_2(original_rsci_idat, aqed_in_if_issue_dup_aif_1_aif_equal_tmp,
      state_orig_issued_sva);
  assign nand_3_nl = ~(mux_5_cse & bmc_v_rsci_idat & duplicate_rsci_idat & (~ state_dup_issued_sva));
  assign state_dup_in_sva_dfm_1_mx1 = MUX_v_16_2_2(state_in_count_sva, state_dup_in_sva,
      nand_3_nl);
  assign nl_aqed_out_if_if_2_acc_nl = ({1'b1 , state_dup_in_sva_dfm_1_mx1}) + conv_u2u_16_17(~
      state_out_count_sva) + 17'b00000000000000001;
  assign aqed_out_if_if_2_acc_nl = nl_aqed_out_if_if_2_acc_nl[16:0];
  assign aqed_out_if_if_2_acc_itm_16_1 = readslicef_17_1_16((aqed_out_if_if_2_acc_nl));
  assign aqed_in_if_aqed_in_if_or_2_nl = state_orig_issued_sva | aqed_in_if_issue_orig_land_lpi_1_dfm_1;
  assign state_orig_issued_sva_dfm_1_mx0 = MUX_s_1_2_2(state_orig_issued_sva, (aqed_in_if_aqed_in_if_or_2_nl),
      bmc_v_rsci_idat);
  assign aqed_in_if_issue_orig_land_lpi_1_dfm_1 = (~ state_orig_issued_sva) & original_rsci_idat;
  assign aqed_in_if_issue_dup_aif_1_aif_equal_tmp = bmc_in_rsci_idat == state_orig_sva;
  assign aqed_in_if_aqed_in_if_or_3_nl = state_dup_issued_sva | ((aqed_in_if_issue_orig_land_lpi_1_dfm_1
      | (aqed_in_if_issue_dup_aif_1_aif_equal_tmp & state_orig_issued_sva)) & duplicate_rsci_idat);
  assign state_dup_issued_sva_mx0 = MUX_s_1_2_2(state_dup_issued_sva, (aqed_in_if_aqed_in_if_or_3_nl),
      bmc_v_rsci_idat);
  assign aqed_out_if_aqed_out_if_and_1_tmp = acc_out_rdy_rsci_idat & acc_out_v_rsci_idat;
  assign and_nl = duplicate_rsci_idat & mux_3_cse;
  assign mux_1_itm = MUX_s_1_2_2((and_nl), or_15_cse, state_dup_issued_sva);
  assign and_dcpl_10 = bmc_v_rsci_idat & clk_en;
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_out_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & (~((mux_1_itm & aqed_out_if_aif_4_equal_tmp) | aqed_out_if_if_2_acc_itm_16_1
        | state_qed_done_sva)) & or_15_cse & aqed_out_if_aqed_out_if_and_1_tmp &
        aqed_out_if_aif_1_equal_tmp ) begin
      state_orig_out_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_out_count_sva <= 16'b0000000000000000;
      state_qed_done_sva <= 1'b0;
      reg_state_orig_done_cse <= 1'b0;
    end
    else if ( state_out_count_and_cse ) begin
      state_out_count_sva <= nl_state_out_count_sva[15:0];
      state_qed_done_sva <= state_qed_done_sva | (aqed_out_if_aif_4_equal_tmp & state_dup_issued_sva_mx0
          & state_orig_issued_sva_dfm_1_mx0) | aqed_out_if_if_2_acc_itm_16_1;
      reg_state_orig_done_cse <= (~ (readslicef_17_1_16((aqed_out_if_aelse_acc_nl))))
          & state_orig_issued_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      reg_state_qed_check_cse <= 1'b0;
    end
    else if ( clk_en & (~((mux_4_nl) | (~(aqed_out_if_aif_4_equal_tmp & aqed_out_if_aqed_out_if_and_1_tmp))
        | state_qed_done_sva)) ) begin
      reg_state_qed_check_cse <= acc_out_rsci_idat == (aqed_out_if_mux_2_nl);
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_dup_in_sva <= 16'b1111111111111111;
    end
    else if ( mux_5_cse & (~ state_dup_issued_sva) & duplicate_rsci_idat & bmc_v_rsci_idat
        & clk_en ) begin
      state_dup_in_sva <= state_dup_in_sva_dfm_1_mx1;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_in_count_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & (~ mux_1_itm) & bmc_v_rsci_idat ) begin
      state_in_count_sva <= nl_state_in_count_sva[15:0];
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_in_sva <= 16'b0000000000000000;
    end
    else if ( and_9_cse & (~ state_orig_issued_sva) & clk_en ) begin
      state_orig_in_sva <= state_orig_in_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & or_15_cse & (~ duplicate_rsci_idat) & (~ state_dup_issued_sva)
        & (~ state_orig_issued_sva) ) begin
      state_orig_sva <= bmc_in_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_issued_sva <= 1'b0;
      state_dup_issued_sva <= 1'b0;
    end
    else if ( and_dcpl_10 ) begin
      state_orig_issued_sva <= state_orig_issued_sva_dfm_1_mx0;
      state_dup_issued_sva <= state_dup_issued_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      return_aqed_out_v_rsci_idat <= 1'b0;
      return_aqed_out_rsci_idat <= 16'b0000000000000000;
    end
    else if ( clk_en ) begin
      return_aqed_out_v_rsci_idat <= bmc_v_rsci_idat;
      return_aqed_out_rsci_idat <= bmc_in_rsci_idat;
    end
  end
  assign nl_state_out_count_sva  = state_out_count_sva + 16'b0000000000000001;
  assign nl_aqed_out_if_aelse_acc_nl = ({1'b1 , state_out_count_sva}) + conv_u2u_16_17(~
      state_orig_in_sva_dfm_1_mx0) + 17'b00000000000000001;
  assign aqed_out_if_aelse_acc_nl = nl_aqed_out_if_aelse_acc_nl[16:0];
  assign aqed_out_if_if_aqed_out_if_if_and_1_nl = (~ state_qed_done_sva) & aqed_out_if_aif_1_equal_tmp
      & state_orig_issued_sva_dfm_1_mx0;
  assign aqed_out_if_mux_2_nl = MUX_v_16_2_2(state_orig_out_sva, acc_out_rsci_idat,
      aqed_out_if_if_aqed_out_if_if_and_1_nl);
  assign nand_1_nl = ~(duplicate_rsci_idat & mux_3_cse);
  assign nor_4_nl = ~(state_orig_issued_sva | and_9_cse);
  assign mux_4_nl = MUX_s_1_2_2((nand_1_nl), (nor_4_nl), state_dup_issued_sva);
  assign nl_state_in_count_sva  = state_in_count_sva + 16'b0000000000000001;

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    aqed_top
// ------------------------------------------------------------------


module aqed_top (
  clk, clk_en, reset, bmc_in_rsc_dat, bmc_v_rsc_dat, original_rsc_dat, duplicate_rsc_dat,
      acc_out_rsc_dat, acc_out_v_rsc_dat, acc_out_rdy_rsc_dat, return_aqed_out_rsc_dat,
      return_aqed_out_v_rsc_dat, return_qed_done_rsc_dat, return_qed_check_rsc_dat,
      return_orig_issued_rsc_dat, return_orig_done_rsc_dat
);
  input clk;
  input clk_en;
  input reset;
  input [15:0] bmc_in_rsc_dat;
  input bmc_v_rsc_dat;
  input original_rsc_dat;
  input duplicate_rsc_dat;
  input [15:0] acc_out_rsc_dat;
  input acc_out_v_rsc_dat;
  input acc_out_rdy_rsc_dat;
  output [15:0] return_aqed_out_rsc_dat;
  output return_aqed_out_v_rsc_dat;
  output return_qed_done_rsc_dat;
  output return_qed_check_rsc_dat;
  output return_orig_issued_rsc_dat;
  output return_orig_done_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  aqed_top_core aqed_top_core_inst (
      .clk(clk),
      .clk_en(clk_en),
      .reset(reset),
      .bmc_in_rsc_dat(bmc_in_rsc_dat),
      .bmc_v_rsc_dat(bmc_v_rsc_dat),
      .original_rsc_dat(original_rsc_dat),
      .duplicate_rsc_dat(duplicate_rsc_dat),
      .acc_out_rsc_dat(acc_out_rsc_dat),
      .acc_out_v_rsc_dat(acc_out_v_rsc_dat),
      .acc_out_rdy_rsc_dat(acc_out_rdy_rsc_dat),
      .return_aqed_out_rsc_dat(return_aqed_out_rsc_dat),
      .return_aqed_out_v_rsc_dat(return_aqed_out_v_rsc_dat),
      .return_qed_done_rsc_dat(return_qed_done_rsc_dat),
      .return_qed_check_rsc_dat(return_qed_check_rsc_dat),
      .return_orig_issued_rsc_dat(return_orig_issued_rsc_dat),
      .return_orig_done_rsc_dat(return_orig_done_rsc_dat)
    );
endmodule



