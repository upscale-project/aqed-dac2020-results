
//------> /hd/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /hd/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   saranyuc@rsg20.stanford.edu
//  Generated date: Sun Mar 29 00:17:46 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    aqed_top_core
// ------------------------------------------------------------------


module aqed_top_core (
  clk, clk_en, reset, bmc_in_rsc_dat, bmc_v_rsc_dat, original_rsc_dat, duplicate_rsc_dat,
      full_rsc_dat, empty_rsc_dat, acc_out_rsc_dat, acc_out_v_rsc_dat, return_aqed_out_rsc_dat,
      return_aqed_out_v_rsc_dat, return_qed_done_rsc_dat, return_qed_check_rsc_dat
);
  input clk;
  input clk_en;
  input reset;
  input [15:0] bmc_in_rsc_dat;
  input bmc_v_rsc_dat;
  input original_rsc_dat;
  input duplicate_rsc_dat;
  input full_rsc_dat;
  input empty_rsc_dat;
  input [15:0] acc_out_rsc_dat;
  input acc_out_v_rsc_dat;
  output [15:0] return_aqed_out_rsc_dat;
  output return_aqed_out_v_rsc_dat;
  output return_qed_done_rsc_dat;
  output return_qed_check_rsc_dat;


  // Interconnect Declarations
  wire [15:0] bmc_in_rsci_idat;
  wire bmc_v_rsci_idat;
  wire original_rsci_idat;
  wire duplicate_rsci_idat;
  wire full_rsci_idat;
  wire empty_rsci_idat;
  wire [15:0] acc_out_rsci_idat;
  wire acc_out_v_rsci_idat;
  reg [15:0] return_aqed_out_rsci_idat;
  reg return_aqed_out_v_rsci_idat;
  reg return_qed_done_rsci_idat;
  reg return_qed_check_rsci_idat;
  wire or_dcpl_2;
  wire not_tmp_7;
  reg state_dup_done_sva;
  reg state_orig_done_sva;
  reg [15:0] state_orig_sva;
  reg state_orig_issued_sva;
  wire [15:0] z_out;
  wire [16:0] nl_z_out;
  reg [15:0] state_orig_in_sva;
  reg [15:0] state_orig_out_sva;
  reg [15:0] state_dup_out_sva;
  reg [15:0] state_dup_in_sva;
  reg [15:0] state_in_count_sva;
  wire [16:0] nl_state_in_count_sva;
  reg [15:0] state_out_count_sva;
  wire [16:0] nl_state_out_count_sva;
  wire [15:0] state_dup_in_sva_dfm_1_mx0;
  wire [15:0] state_orig_in_sva_dfm_1_mx0;
  wire [15:0] state_dup_out_sva_dfm_1_mx0;
  wire [15:0] state_orig_out_sva_dfm_1_mx0;
  wire state_dup_done_sva_mx0;
  wire state_orig_done_sva_mx0;
  wire equal_tmp;
  wire and_9_cse;
  wire and_19_cse;
  wire aqed_out_if_if_1_acc_itm_16;
  wire aqed_out_if_if_acc_itm_16;

  wire[0:0] or_4_nl;
  wire[0:0] or_6_nl;
  wire[0:0] or_8_nl;
  wire[16:0] aqed_out_if_if_1_acc_nl;
  wire[18:0] nl_aqed_out_if_if_1_acc_nl;
  wire[0:0] or_10_nl;
  wire[16:0] aqed_out_if_if_acc_nl;
  wire[18:0] nl_aqed_out_if_if_acc_nl;
  wire[0:0] aqed_out_if_aqed_out_if_or_2_nl;
  wire[0:0] aqed_out_if_aqed_out_if_or_3_nl;
  wire[0:0] aqed_in_if_if_1_mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd16)) bmc_in_rsci (
      .dat(bmc_in_rsc_dat),
      .idat(bmc_in_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd1)) bmc_v_rsci (
      .dat(bmc_v_rsc_dat),
      .idat(bmc_v_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd1)) original_rsci (
      .dat(original_rsc_dat),
      .idat(original_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd1)) duplicate_rsci (
      .dat(duplicate_rsc_dat),
      .idat(duplicate_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd1)) full_rsci (
      .dat(full_rsc_dat),
      .idat(full_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd1)) empty_rsci (
      .dat(empty_rsc_dat),
      .idat(empty_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd16)) acc_out_rsci (
      .dat(acc_out_rsc_dat),
      .idat(acc_out_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd1)) acc_out_v_rsci (
      .dat(acc_out_v_rsc_dat),
      .idat(acc_out_v_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd9),
  .width(32'sd16)) return_aqed_out_rsci (
      .idat(return_aqed_out_rsci_idat),
      .dat(return_aqed_out_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd10),
  .width(32'sd1)) return_aqed_out_v_rsci (
      .idat(return_aqed_out_v_rsci_idat),
      .dat(return_aqed_out_v_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd11),
  .width(32'sd1)) return_qed_done_rsci (
      .idat(return_qed_done_rsci_idat),
      .dat(return_qed_done_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd12),
  .width(32'sd1)) return_qed_check_rsci (
      .idat(return_qed_check_rsci_idat),
      .dat(return_qed_check_rsc_dat)
    );
  assign and_9_cse = (~ state_orig_issued_sva) & original_rsci_idat & (~ full_rsci_idat)
      & clk_en & bmc_v_rsci_idat;
  assign and_19_cse = acc_out_v_rsci_idat & (~ empty_rsci_idat) & clk_en;
  assign equal_tmp = bmc_in_rsci_idat == state_orig_sva;
  assign or_4_nl = or_dcpl_2 | (~ state_orig_issued_sva) | (~(duplicate_rsci_idat
      & equal_tmp));
  assign state_dup_in_sva_dfm_1_mx0 = MUX_v_16_2_2(z_out, state_dup_in_sva, or_4_nl);
  assign or_6_nl = or_dcpl_2 | (~ original_rsci_idat) | state_orig_issued_sva;
  assign state_orig_in_sva_dfm_1_mx0 = MUX_v_16_2_2(z_out, state_orig_in_sva, or_6_nl);
  assign or_8_nl = not_tmp_7 | aqed_out_if_if_1_acc_itm_16 | state_dup_done_sva;
  assign state_dup_out_sva_dfm_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_dup_out_sva,
      or_8_nl);
  assign nl_aqed_out_if_if_1_acc_nl = ({1'b1 , state_out_count_sva}) + conv_u2u_16_17(~
      state_dup_in_sva_dfm_1_mx0) + 17'b00000000000000001;
  assign aqed_out_if_if_1_acc_nl = nl_aqed_out_if_if_1_acc_nl[16:0];
  assign aqed_out_if_if_1_acc_itm_16 = readslicef_17_1_16((aqed_out_if_if_1_acc_nl));
  assign or_10_nl = not_tmp_7 | aqed_out_if_if_acc_itm_16 | state_orig_done_sva;
  assign state_orig_out_sva_dfm_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_orig_out_sva,
      or_10_nl);
  assign nl_aqed_out_if_if_acc_nl = ({1'b1 , state_out_count_sva}) + conv_u2u_16_17(~
      state_orig_in_sva_dfm_1_mx0) + 17'b00000000000000001;
  assign aqed_out_if_if_acc_nl = nl_aqed_out_if_if_acc_nl[16:0];
  assign aqed_out_if_if_acc_itm_16 = readslicef_17_1_16((aqed_out_if_if_acc_nl));
  assign aqed_out_if_aqed_out_if_or_2_nl = state_dup_done_sva | (~ aqed_out_if_if_1_acc_itm_16);
  assign state_dup_done_sva_mx0 = MUX_s_1_2_2((aqed_out_if_aqed_out_if_or_2_nl),
      state_dup_done_sva, not_tmp_7);
  assign aqed_out_if_aqed_out_if_or_3_nl = state_orig_done_sva | (~ aqed_out_if_if_acc_itm_16);
  assign state_orig_done_sva_mx0 = MUX_s_1_2_2((aqed_out_if_aqed_out_if_or_3_nl),
      state_orig_done_sva, not_tmp_7);
  assign or_dcpl_2 = (~ bmc_v_rsci_idat) | full_rsci_idat;
  assign not_tmp_7 = ~((~ empty_rsci_idat) & acc_out_v_rsci_idat);
  always @(posedge clk) begin
    if ( reset ) begin
      state_dup_in_sva <= 16'b1111111111111111;
    end
    else if ( equal_tmp & duplicate_rsci_idat & state_orig_issued_sva & (~ full_rsci_idat)
        & clk_en & bmc_v_rsci_idat ) begin
      state_dup_in_sva <= state_dup_in_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_in_sva <= 16'b1111111111111111;
      state_orig_sva <= 16'b0000000000000000;
    end
    else if ( and_9_cse ) begin
      state_orig_in_sva <= state_orig_in_sva_dfm_1_mx0;
      state_orig_sva <= bmc_in_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_in_count_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & (~ or_dcpl_2) ) begin
      state_in_count_sva <= nl_state_in_count_sva[15:0];
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_issued_sva <= 1'b0;
      return_qed_check_rsci_idat <= 1'b0;
      return_qed_done_rsci_idat <= 1'b0;
      return_aqed_out_v_rsci_idat <= 1'b0;
      return_aqed_out_rsci_idat <= 16'b0000000000000000;
    end
    else if ( clk_en ) begin
      state_orig_issued_sva <= state_orig_issued_sva | (original_rsci_idat & (~(full_rsci_idat
          | (~ bmc_v_rsci_idat))));
      return_qed_check_rsci_idat <= state_orig_out_sva_dfm_1_mx0 == state_dup_out_sva_dfm_1_mx0;
      return_qed_done_rsci_idat <= state_dup_done_sva_mx0 & state_orig_done_sva_mx0;
      return_aqed_out_v_rsci_idat <= bmc_v_rsci_idat;
      return_aqed_out_rsci_idat <= bmc_in_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_dup_out_sva <= 16'b0000000000000000;
    end
    else if ( (~(state_dup_done_sva | aqed_out_if_if_1_acc_itm_16)) & acc_out_v_rsci_idat
        & clk_en & (~ empty_rsci_idat) ) begin
      state_dup_out_sva <= state_dup_out_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_out_sva <= 16'b0000000000000000;
    end
    else if ( (~(state_orig_done_sva | aqed_out_if_if_acc_itm_16)) & acc_out_v_rsci_idat
        & clk_en & (~ empty_rsci_idat) ) begin
      state_orig_out_sva <= state_orig_out_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_dup_done_sva <= 1'b0;
      state_orig_done_sva <= 1'b0;
    end
    else if ( and_19_cse ) begin
      state_dup_done_sva <= state_dup_done_sva_mx0;
      state_orig_done_sva <= state_orig_done_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_out_count_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & (~ not_tmp_7) ) begin
      state_out_count_sva <= nl_state_out_count_sva[15:0];
    end
  end
  assign nl_state_in_count_sva  = state_in_count_sva + 16'b0000000000000001;
  assign nl_state_out_count_sva  = state_out_count_sva + 16'b0000000000000001;
  assign aqed_in_if_if_1_mux_1_nl = MUX_s_1_2_2((~ original_rsci_idat), (~ duplicate_rsci_idat),
      state_orig_issued_sva);
  assign nl_z_out = state_in_count_sva + conv_s2u_1_16(aqed_in_if_if_1_mux_1_nl);
  assign z_out = nl_z_out[15:0];

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [15:0] conv_s2u_1_16 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_16 = {{15{vector[0]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    aqed_top
// ------------------------------------------------------------------


module aqed_top (
  clk, clk_en, reset, bmc_in_rsc_dat, bmc_v_rsc_dat, original_rsc_dat, duplicate_rsc_dat,
      full_rsc_dat, empty_rsc_dat, acc_out_rsc_dat, acc_out_v_rsc_dat, return_aqed_out_rsc_dat,
      return_aqed_out_v_rsc_dat, return_qed_done_rsc_dat, return_qed_check_rsc_dat
);
  input clk;
  input clk_en;
  input reset;
  input [15:0] bmc_in_rsc_dat;
  input bmc_v_rsc_dat;
  input original_rsc_dat;
  input duplicate_rsc_dat;
  input full_rsc_dat;
  input empty_rsc_dat;
  input [15:0] acc_out_rsc_dat;
  input acc_out_v_rsc_dat;
  output [15:0] return_aqed_out_rsc_dat;
  output return_aqed_out_v_rsc_dat;
  output return_qed_done_rsc_dat;
  output return_qed_check_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  aqed_top_core aqed_top_core_inst (
      .clk(clk),
      .clk_en(clk_en),
      .reset(reset),
      .bmc_in_rsc_dat(bmc_in_rsc_dat),
      .bmc_v_rsc_dat(bmc_v_rsc_dat),
      .original_rsc_dat(original_rsc_dat),
      .duplicate_rsc_dat(duplicate_rsc_dat),
      .full_rsc_dat(full_rsc_dat),
      .empty_rsc_dat(empty_rsc_dat),
      .acc_out_rsc_dat(acc_out_rsc_dat),
      .acc_out_v_rsc_dat(acc_out_v_rsc_dat),
      .return_aqed_out_rsc_dat(return_aqed_out_rsc_dat),
      .return_aqed_out_v_rsc_dat(return_aqed_out_v_rsc_dat),
      .return_qed_done_rsc_dat(return_qed_done_rsc_dat),
      .return_qed_check_rsc_dat(return_qed_check_rsc_dat)
    );
endmodule



