
//------> /hd/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /hd/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   saranyuc@rsg20.stanford.edu
//  Generated date: Fri Apr  3 19:52:37 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    aqed_top_core
// ------------------------------------------------------------------


module aqed_top_core (
  clk, clk_en, reset, bmc_in_rsc_dat, bmc_v_rsc_dat, original_rsc_dat, duplicate_rsc_dat,
      acc_out_rsc_dat, acc_out_v_rsc_dat, acc_out_rdy_rsc_dat, return_aqed_out_rsc_dat,
      return_aqed_out_v_rsc_dat, return_qed_done_rsc_dat, return_qed_check_rsc_dat,
      return_orig_issued_rsc_dat, return_orig_done_rsc_dat
);
  input clk;
  input clk_en;
  input reset;
  input [15:0] bmc_in_rsc_dat;
  input bmc_v_rsc_dat;
  input original_rsc_dat;
  input duplicate_rsc_dat;
  input [15:0] acc_out_rsc_dat;
  input acc_out_v_rsc_dat;
  input acc_out_rdy_rsc_dat;
  output [15:0] return_aqed_out_rsc_dat;
  output return_aqed_out_v_rsc_dat;
  output return_qed_done_rsc_dat;
  output return_qed_check_rsc_dat;
  output return_orig_issued_rsc_dat;
  output return_orig_done_rsc_dat;


  // Interconnect Declarations
  wire [15:0] bmc_in_rsci_idat;
  wire bmc_v_rsci_idat;
  wire original_rsci_idat;
  wire duplicate_rsci_idat;
  wire [15:0] acc_out_rsci_idat;
  wire acc_out_v_rsci_idat;
  wire acc_out_rdy_rsci_idat;
  reg [15:0] return_aqed_out_rsci_idat;
  reg return_aqed_out_v_rsci_idat;
  wire aqed_out_if_aqed_out_if_and_1_tmp;
  wire aqed_in_if_issue_dup_aif_1_aif_equal_tmp;
  wire and_dcpl;
  wire or_dcpl_4;
  wire or_dcpl_5;
  wire or_dcpl_6;
  wire or_dcpl_7;
  wire or_dcpl_8;
  wire or_dcpl_10;
  wire or_dcpl_12;
  wire or_dcpl_13;
  wire or_dcpl_16;
  wire or_dcpl_17;
  wire or_dcpl_20;
  wire or_dcpl_21;
  wire or_dcpl_24;
  wire or_dcpl_25;
  wire or_dcpl_27;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_39;
  wire or_dcpl_42;
  wire or_dcpl_45;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire or_dcpl_60;
  wire or_dcpl_63;
  wire or_dcpl_66;
  wire or_dcpl_77;
  wire or_dcpl_78;
  wire or_dcpl_81;
  wire or_dcpl_84;
  wire or_dcpl_87;
  wire or_dcpl_98;
  wire or_dcpl_99;
  wire or_dcpl_101;
  wire or_dcpl_109;
  wire or_dcpl_110;
  wire or_dcpl_112;
  wire or_dcpl_168;
  wire or_dcpl_169;
  wire or_dcpl_171;
  wire or_dcpl_172;
  wire or_dcpl_174;
  wire or_dcpl_176;
  wire or_dcpl_190;
  wire or_dcpl_192;
  wire or_dcpl_194;
  wire or_dcpl_196;
  reg state_qed_done_sva;
  wire state_dup_issued_sva_mx0;
  wire state_orig_issued_sva_mx0;
  wire aqed_in_if_issue_orig_land_lpi_1_dfm_1;
  reg state_orig_issued_sva;
  reg state_dup_issued_sva;
  reg [15:0] state_out_count_sva;
  wire [16:0] nl_state_out_count_sva;
  reg reg_state_orig_done_cse;
  reg reg_state_qed_check_cse;
  wire and_9_cse;
  wire state_out_count_and_cse;
  wire mux_6_cse;
  reg [15:0] state_orig_in_sva;
  reg [15:0] state_dup_in_sva;
  reg [15:0] state_in_count_sva;
  wire [16:0] nl_state_in_count_sva;
  reg [15:0] state_output_63_sva;
  reg [15:0] state_output_64_sva;
  reg [15:0] state_output_62_sva;
  reg [15:0] state_output_65_sva;
  reg [15:0] state_output_61_sva;
  reg [15:0] state_output_66_sva;
  reg [15:0] state_output_60_sva;
  reg [15:0] state_output_67_sva;
  reg [15:0] state_output_59_sva;
  reg [15:0] state_output_68_sva;
  reg [15:0] state_output_58_sva;
  reg [15:0] state_output_69_sva;
  reg [15:0] state_output_57_sva;
  reg [15:0] state_output_70_sva;
  reg [15:0] state_output_56_sva;
  reg [15:0] state_output_71_sva;
  reg [15:0] state_output_55_sva;
  reg [15:0] state_output_72_sva;
  reg [15:0] state_output_54_sva;
  reg [15:0] state_output_73_sva;
  reg [15:0] state_output_53_sva;
  reg [15:0] state_output_74_sva;
  reg [15:0] state_output_52_sva;
  reg [15:0] state_output_75_sva;
  reg [15:0] state_output_51_sva;
  reg [15:0] state_output_76_sva;
  reg [15:0] state_output_50_sva;
  reg [15:0] state_output_77_sva;
  reg [15:0] state_output_49_sva;
  reg [15:0] state_output_78_sva;
  reg [15:0] state_output_48_sva;
  reg [15:0] state_output_79_sva;
  reg [15:0] state_output_47_sva;
  reg [15:0] state_output_80_sva;
  reg [15:0] state_output_46_sva;
  reg [15:0] state_output_81_sva;
  reg [15:0] state_output_45_sva;
  reg [15:0] state_output_82_sva;
  reg [15:0] state_output_44_sva;
  reg [15:0] state_output_83_sva;
  reg [15:0] state_output_43_sva;
  reg [15:0] state_output_84_sva;
  reg [15:0] state_output_42_sva;
  reg [15:0] state_output_85_sva;
  reg [15:0] state_output_41_sva;
  reg [15:0] state_output_86_sva;
  reg [15:0] state_output_40_sva;
  reg [15:0] state_output_87_sva;
  reg [15:0] state_output_39_sva;
  reg [15:0] state_output_88_sva;
  reg [15:0] state_output_38_sva;
  reg [15:0] state_output_89_sva;
  reg [15:0] state_output_37_sva;
  reg [15:0] state_output_90_sva;
  reg [15:0] state_output_36_sva;
  reg [15:0] state_output_91_sva;
  reg [15:0] state_output_35_sva;
  reg [15:0] state_output_92_sva;
  reg [15:0] state_output_34_sva;
  reg [15:0] state_output_93_sva;
  reg [15:0] state_output_33_sva;
  reg [15:0] state_output_94_sva;
  reg [15:0] state_output_32_sva;
  reg [15:0] state_output_95_sva;
  reg [15:0] state_output_31_sva;
  reg [15:0] state_output_96_sva;
  reg [15:0] state_output_30_sva;
  reg [15:0] state_output_97_sva;
  reg [15:0] state_output_29_sva;
  reg [15:0] state_output_98_sva;
  reg [15:0] state_output_28_sva;
  reg [15:0] state_output_99_sva;
  reg [15:0] state_output_27_sva;
  reg [15:0] state_output_100_sva;
  reg [15:0] state_output_26_sva;
  reg [15:0] state_output_101_sva;
  reg [15:0] state_output_25_sva;
  reg [15:0] state_output_102_sva;
  reg [15:0] state_output_24_sva;
  reg [15:0] state_output_103_sva;
  reg [15:0] state_output_23_sva;
  reg [15:0] state_output_104_sva;
  reg [15:0] state_output_22_sva;
  reg [15:0] state_output_105_sva;
  reg [15:0] state_output_21_sva;
  reg [15:0] state_output_106_sva;
  reg [15:0] state_output_20_sva;
  reg [15:0] state_output_107_sva;
  reg [15:0] state_output_19_sva;
  reg [15:0] state_output_108_sva;
  reg [15:0] state_output_18_sva;
  reg [15:0] state_output_109_sva;
  reg [15:0] state_output_17_sva;
  reg [15:0] state_output_110_sva;
  reg [15:0] state_output_16_sva;
  reg [15:0] state_output_111_sva;
  reg [15:0] state_output_15_sva;
  reg [15:0] state_output_112_sva;
  reg [15:0] state_output_14_sva;
  reg [15:0] state_output_113_sva;
  reg [15:0] state_output_13_sva;
  reg [15:0] state_output_114_sva;
  reg [15:0] state_output_12_sva;
  reg [15:0] state_output_115_sva;
  reg [15:0] state_output_11_sva;
  reg [15:0] state_output_116_sva;
  reg [15:0] state_output_10_sva;
  reg [15:0] state_output_117_sva;
  reg [15:0] state_output_9_sva;
  reg [15:0] state_output_118_sva;
  reg [15:0] state_output_8_sva;
  reg [15:0] state_output_119_sva;
  reg [15:0] state_output_7_sva;
  reg [15:0] state_output_120_sva;
  reg [15:0] state_output_6_sva;
  reg [15:0] state_output_121_sva;
  reg [15:0] state_output_5_sva;
  reg [15:0] state_output_122_sva;
  reg [15:0] state_output_4_sva;
  reg [15:0] state_output_123_sva;
  reg [15:0] state_output_3_sva;
  reg [15:0] state_output_124_sva;
  reg [15:0] state_output_2_sva;
  reg [15:0] state_output_125_sva;
  reg [15:0] state_output_1_sva;
  reg [15:0] state_output_126_sva;
  reg [15:0] state_output_0_sva;
  reg [15:0] state_output_127_sva;
  reg state_orig_idx_sva;
  reg state_dup_idx_sva;
  wire [15:0] state_orig_in_sva_dfm_1_mx0;
  wire [15:0] state_output_0_sva_1_mx0;
  wire [15:0] state_output_1_sva_1_mx0;
  wire [15:0] state_output_2_sva_1_mx0;
  wire [15:0] state_output_3_sva_1_mx0;
  wire [15:0] state_output_4_sva_1_mx0;
  wire [15:0] state_output_5_sva_1_mx0;
  wire [15:0] state_output_6_sva_1_mx0;
  wire [15:0] state_output_7_sva_1_mx0;
  wire [15:0] state_output_8_sva_1_mx0;
  wire [15:0] state_output_9_sva_1_mx0;
  wire [15:0] state_output_10_sva_1_mx0;
  wire [15:0] state_output_11_sva_1_mx0;
  wire [15:0] state_output_12_sva_1_mx0;
  wire [15:0] state_output_13_sva_1_mx0;
  wire [15:0] state_output_14_sva_1_mx0;
  wire [15:0] state_output_15_sva_1_mx0;
  wire [15:0] state_output_16_sva_1_mx0;
  wire [15:0] state_output_17_sva_1_mx0;
  wire [15:0] state_output_18_sva_1_mx0;
  wire [15:0] state_output_19_sva_1_mx0;
  wire [15:0] state_output_20_sva_1_mx0;
  wire [15:0] state_output_21_sva_1_mx0;
  wire [15:0] state_output_22_sva_1_mx0;
  wire [15:0] state_output_23_sva_1_mx0;
  wire [15:0] state_output_24_sva_1_mx0;
  wire [15:0] state_output_25_sva_1_mx0;
  wire [15:0] state_output_26_sva_1_mx0;
  wire [15:0] state_output_27_sva_1_mx0;
  wire [15:0] state_output_28_sva_1_mx0;
  wire [15:0] state_output_29_sva_1_mx0;
  wire [15:0] state_output_30_sva_1_mx0;
  wire [15:0] state_output_31_sva_1_mx0;
  wire [15:0] state_output_32_sva_1_mx0;
  wire [15:0] state_output_33_sva_1_mx0;
  wire [15:0] state_output_34_sva_1_mx0;
  wire [15:0] state_output_35_sva_1_mx0;
  wire [15:0] state_output_36_sva_1_mx0;
  wire [15:0] state_output_37_sva_1_mx0;
  wire [15:0] state_output_38_sva_1_mx0;
  wire [15:0] state_output_39_sva_1_mx0;
  wire [15:0] state_output_40_sva_1_mx0;
  wire [15:0] state_output_41_sva_1_mx0;
  wire [15:0] state_output_42_sva_1_mx0;
  wire [15:0] state_output_43_sva_1_mx0;
  wire [15:0] state_output_44_sva_1_mx0;
  wire [15:0] state_output_45_sva_1_mx0;
  wire [15:0] state_output_46_sva_1_mx0;
  wire [15:0] state_output_47_sva_1_mx0;
  wire [15:0] state_output_48_sva_1_mx0;
  wire [15:0] state_output_49_sva_1_mx0;
  wire [15:0] state_output_50_sva_1_mx0;
  wire [15:0] state_output_51_sva_1_mx0;
  wire [15:0] state_output_52_sva_1_mx0;
  wire [15:0] state_output_53_sva_1_mx0;
  wire [15:0] state_output_54_sva_1_mx0;
  wire [15:0] state_output_55_sva_1_mx0;
  wire [15:0] state_output_56_sva_1_mx0;
  wire [15:0] state_output_57_sva_1_mx0;
  wire [15:0] state_output_58_sva_1_mx0;
  wire [15:0] state_output_59_sva_1_mx0;
  wire [15:0] state_output_60_sva_1_mx0;
  wire [15:0] state_output_61_sva_1_mx0;
  wire [15:0] state_output_62_sva_1_mx0;
  wire [15:0] state_output_63_sva_1_mx0;
  wire [15:0] state_output_64_sva_1_mx0;
  wire [15:0] state_output_65_sva_1_mx0;
  wire [15:0] state_output_66_sva_1_mx0;
  wire [15:0] state_output_67_sva_1_mx0;
  wire [15:0] state_output_68_sva_1_mx0;
  wire [15:0] state_output_69_sva_1_mx0;
  wire [15:0] state_output_70_sva_1_mx0;
  wire [15:0] state_output_71_sva_1_mx0;
  wire [15:0] state_output_72_sva_1_mx0;
  wire [15:0] state_output_73_sva_1_mx0;
  wire [15:0] state_output_74_sva_1_mx0;
  wire [15:0] state_output_75_sva_1_mx0;
  wire [15:0] state_output_76_sva_1_mx0;
  wire [15:0] state_output_77_sva_1_mx0;
  wire [15:0] state_output_78_sva_1_mx0;
  wire [15:0] state_output_79_sva_1_mx0;
  wire [15:0] state_output_80_sva_1_mx0;
  wire [15:0] state_output_81_sva_1_mx0;
  wire [15:0] state_output_82_sva_1_mx0;
  wire [15:0] state_output_83_sva_1_mx0;
  wire [15:0] state_output_84_sva_1_mx0;
  wire [15:0] state_output_85_sva_1_mx0;
  wire [15:0] state_output_86_sva_1_mx0;
  wire [15:0] state_output_87_sva_1_mx0;
  wire [15:0] state_output_88_sva_1_mx0;
  wire [15:0] state_output_89_sva_1_mx0;
  wire [15:0] state_output_90_sva_1_mx0;
  wire [15:0] state_output_91_sva_1_mx0;
  wire [15:0] state_output_92_sva_1_mx0;
  wire [15:0] state_output_93_sva_1_mx0;
  wire [15:0] state_output_94_sva_1_mx0;
  wire [15:0] state_output_95_sva_1_mx0;
  wire [15:0] state_output_96_sva_1_mx0;
  wire [15:0] state_output_97_sva_1_mx0;
  wire [15:0] state_output_98_sva_1_mx0;
  wire [15:0] state_output_99_sva_1_mx0;
  wire [15:0] state_output_100_sva_1_mx0;
  wire [15:0] state_output_101_sva_1_mx0;
  wire [15:0] state_output_102_sva_1_mx0;
  wire [15:0] state_output_103_sva_1_mx0;
  wire [15:0] state_output_104_sva_1_mx0;
  wire [15:0] state_output_105_sva_1_mx0;
  wire [15:0] state_output_106_sva_1_mx0;
  wire [15:0] state_output_107_sva_1_mx0;
  wire [15:0] state_output_108_sva_1_mx0;
  wire [15:0] state_output_109_sva_1_mx0;
  wire [15:0] state_output_110_sva_1_mx0;
  wire [15:0] state_output_111_sva_1_mx0;
  wire [15:0] state_output_112_sva_1_mx0;
  wire [15:0] state_output_113_sva_1_mx0;
  wire [15:0] state_output_114_sva_1_mx0;
  wire [15:0] state_output_115_sva_1_mx0;
  wire [15:0] state_output_116_sva_1_mx0;
  wire [15:0] state_output_117_sva_1_mx0;
  wire [15:0] state_output_118_sva_1_mx0;
  wire [15:0] state_output_119_sva_1_mx0;
  wire [15:0] state_output_120_sva_1_mx0;
  wire [15:0] state_output_121_sva_1_mx0;
  wire [15:0] state_output_122_sva_1_mx0;
  wire [15:0] state_output_123_sva_1_mx0;
  wire [15:0] state_output_124_sva_1_mx0;
  wire [15:0] state_output_125_sva_1_mx0;
  wire [15:0] state_output_126_sva_1_mx0;
  wire [15:0] state_output_127_sva_1_mx0;
  wire state_orig_idx_sva_dfm_1_mx0;
  wire [15:0] state_dup_in_sva_dfm_1_mx0;
  wire state_dup_idx_sva_dfm_1_mx0;
  wire aqed_in_if_issue_dup_land_1_lpi_1_dfm_2;
  wire nor_10_rgt;
  wire and_dcpl_23;
  wire aqed_out_if_aelse_2_acc_itm_16;

  wire[0:0] mux_5_nl;
  wire[0:0] and_8_nl;
  wire[0:0] and_11_nl;
  wire[0:0] or_316_nl;
  wire[15:0] aqed_out_if_if_mux_nl;
  wire[6:0] operator_ac_int_16_false_1_false_2_acc_nl;
  wire[7:0] nl_operator_ac_int_16_false_1_false_2_acc_nl;
  wire[15:0] aqed_out_if_if_mux_3_nl;
  wire[6:0] operator_ac_int_16_false_1_false_3_acc_nl;
  wire[7:0] nl_operator_ac_int_16_false_1_false_3_acc_nl;
  wire[0:0] mux_nl;
  wire[16:0] aqed_out_if_aelse_acc_nl;
  wire[18:0] nl_aqed_out_if_aelse_acc_nl;
  wire[0:0] or_17_nl;
  wire[0:0] or_19_nl;
  wire[0:0] or_22_nl;
  wire[0:0] or_23_nl;
  wire[0:0] or_26_nl;
  wire[0:0] or_27_nl;
  wire[0:0] or_30_nl;
  wire[0:0] or_31_nl;
  wire[0:0] or_34_nl;
  wire[0:0] or_36_nl;
  wire[0:0] or_37_nl;
  wire[0:0] or_38_nl;
  wire[0:0] or_39_nl;
  wire[0:0] or_40_nl;
  wire[0:0] or_41_nl;
  wire[0:0] or_42_nl;
  wire[0:0] or_45_nl;
  wire[0:0] or_46_nl;
  wire[0:0] or_48_nl;
  wire[0:0] or_49_nl;
  wire[0:0] or_51_nl;
  wire[0:0] or_52_nl;
  wire[0:0] or_54_nl;
  wire[0:0] or_55_nl;
  wire[0:0] or_56_nl;
  wire[0:0] or_57_nl;
  wire[0:0] or_58_nl;
  wire[0:0] or_59_nl;
  wire[0:0] or_60_nl;
  wire[0:0] or_61_nl;
  wire[0:0] or_62_nl;
  wire[0:0] or_63_nl;
  wire[0:0] or_66_nl;
  wire[0:0] or_67_nl;
  wire[0:0] or_69_nl;
  wire[0:0] or_70_nl;
  wire[0:0] or_72_nl;
  wire[0:0] or_73_nl;
  wire[0:0] or_75_nl;
  wire[0:0] or_76_nl;
  wire[0:0] or_77_nl;
  wire[0:0] or_78_nl;
  wire[0:0] or_79_nl;
  wire[0:0] or_80_nl;
  wire[0:0] or_81_nl;
  wire[0:0] or_82_nl;
  wire[0:0] or_83_nl;
  wire[0:0] or_84_nl;
  wire[0:0] or_87_nl;
  wire[0:0] or_88_nl;
  wire[0:0] or_90_nl;
  wire[0:0] or_91_nl;
  wire[0:0] or_93_nl;
  wire[0:0] or_94_nl;
  wire[0:0] or_96_nl;
  wire[0:0] or_97_nl;
  wire[0:0] or_98_nl;
  wire[0:0] or_99_nl;
  wire[0:0] or_100_nl;
  wire[0:0] or_101_nl;
  wire[0:0] or_102_nl;
  wire[0:0] or_103_nl;
  wire[0:0] or_104_nl;
  wire[0:0] or_105_nl;
  wire[0:0] or_108_nl;
  wire[0:0] or_110_nl;
  wire[0:0] or_111_nl;
  wire[0:0] or_112_nl;
  wire[0:0] or_113_nl;
  wire[0:0] or_114_nl;
  wire[0:0] or_115_nl;
  wire[0:0] or_116_nl;
  wire[0:0] or_119_nl;
  wire[0:0] or_121_nl;
  wire[0:0] or_122_nl;
  wire[0:0] or_123_nl;
  wire[0:0] or_124_nl;
  wire[0:0] or_125_nl;
  wire[0:0] or_126_nl;
  wire[0:0] or_127_nl;
  wire[0:0] or_128_nl;
  wire[0:0] or_129_nl;
  wire[0:0] or_130_nl;
  wire[0:0] or_131_nl;
  wire[0:0] or_132_nl;
  wire[0:0] or_133_nl;
  wire[0:0] or_134_nl;
  wire[0:0] or_135_nl;
  wire[0:0] or_136_nl;
  wire[0:0] or_137_nl;
  wire[0:0] or_138_nl;
  wire[0:0] or_139_nl;
  wire[0:0] or_140_nl;
  wire[0:0] or_141_nl;
  wire[0:0] or_142_nl;
  wire[0:0] or_143_nl;
  wire[0:0] or_144_nl;
  wire[0:0] or_145_nl;
  wire[0:0] or_146_nl;
  wire[0:0] or_147_nl;
  wire[0:0] or_148_nl;
  wire[0:0] or_149_nl;
  wire[0:0] or_150_nl;
  wire[0:0] or_151_nl;
  wire[0:0] or_152_nl;
  wire[0:0] or_153_nl;
  wire[0:0] or_154_nl;
  wire[0:0] or_155_nl;
  wire[0:0] or_156_nl;
  wire[0:0] or_157_nl;
  wire[0:0] or_158_nl;
  wire[0:0] or_159_nl;
  wire[0:0] or_160_nl;
  wire[0:0] or_161_nl;
  wire[0:0] or_162_nl;
  wire[0:0] or_163_nl;
  wire[0:0] or_164_nl;
  wire[0:0] or_165_nl;
  wire[0:0] or_166_nl;
  wire[0:0] or_167_nl;
  wire[0:0] or_168_nl;
  wire[0:0] or_169_nl;
  wire[0:0] or_170_nl;
  wire[0:0] or_171_nl;
  wire[0:0] or_172_nl;
  wire[0:0] or_173_nl;
  wire[0:0] or_174_nl;
  wire[0:0] or_175_nl;
  wire[0:0] aqed_in_if_mux_7_nl;
  wire[0:0] aqed_in_if_mux_8_nl;
  wire[16:0] aqed_out_if_aelse_2_acc_nl;
  wire[18:0] nl_aqed_out_if_aelse_2_acc_nl;
  wire[0:0] aqed_in_if_aqed_in_if_or_2_nl;
  wire[0:0] aqed_in_if_aqed_in_if_or_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_return_qed_done_rsci_idat;
  assign nl_return_qed_done_rsci_idat = state_qed_done_sva;
  wire [0:0] nl_return_qed_check_rsci_idat;
  assign nl_return_qed_check_rsci_idat = reg_state_qed_check_cse;
  wire [0:0] nl_return_orig_issued_rsci_idat;
  assign nl_return_orig_issued_rsci_idat = state_orig_issued_sva;
  wire [0:0] nl_return_orig_done_rsci_idat;
  assign nl_return_orig_done_rsci_idat = reg_state_orig_done_cse;
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd16)) bmc_in_rsci (
      .dat(bmc_in_rsc_dat),
      .idat(bmc_in_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd1)) bmc_v_rsci (
      .dat(bmc_v_rsc_dat),
      .idat(bmc_v_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd1)) original_rsci (
      .dat(original_rsc_dat),
      .idat(original_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd1)) duplicate_rsci (
      .dat(duplicate_rsc_dat),
      .idat(duplicate_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd16)) acc_out_rsci (
      .dat(acc_out_rsc_dat),
      .idat(acc_out_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd1)) acc_out_v_rsci (
      .dat(acc_out_v_rsc_dat),
      .idat(acc_out_v_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd1)) acc_out_rdy_rsci (
      .dat(acc_out_rdy_rsc_dat),
      .idat(acc_out_rdy_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd8),
  .width(32'sd16)) return_aqed_out_rsci (
      .idat(return_aqed_out_rsci_idat),
      .dat(return_aqed_out_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd9),
  .width(32'sd1)) return_aqed_out_v_rsci (
      .idat(return_aqed_out_v_rsci_idat),
      .dat(return_aqed_out_v_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd10),
  .width(32'sd1)) return_qed_done_rsci (
      .idat(nl_return_qed_done_rsci_idat[0:0]),
      .dat(return_qed_done_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd11),
  .width(32'sd1)) return_qed_check_rsci (
      .idat(nl_return_qed_check_rsci_idat[0:0]),
      .dat(return_qed_check_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd12),
  .width(32'sd1)) return_orig_issued_rsci (
      .idat(nl_return_orig_issued_rsci_idat[0:0]),
      .dat(return_orig_issued_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd13),
  .width(32'sd1)) return_orig_done_rsci (
      .idat(nl_return_orig_done_rsci_idat[0:0]),
      .dat(return_orig_done_rsc_dat)
    );
  assign state_out_count_and_cse = clk_en & aqed_out_if_aqed_out_if_and_1_tmp;
  assign and_8_nl = duplicate_rsci_idat & original_rsci_idat & bmc_v_rsci_idat;
  assign and_11_nl = duplicate_rsci_idat & bmc_v_rsci_idat & aqed_in_if_issue_dup_aif_1_aif_equal_tmp;
  assign mux_5_nl = MUX_s_1_2_2((and_8_nl), (and_11_nl), state_orig_issued_sva);
  assign or_316_nl = state_orig_issued_sva | and_9_cse;
  assign mux_6_cse = MUX_s_1_2_2((mux_5_nl), (or_316_nl), state_dup_issued_sva);
  assign nor_10_rgt = ~(duplicate_rsci_idat | state_orig_issued_sva | state_dup_issued_sva);
  assign state_orig_in_sva_dfm_1_mx0 = MUX_v_16_2_2(state_in_count_sva, state_orig_in_sva,
      state_orig_issued_sva);
  assign or_17_nl = or_dcpl_8 | or_dcpl_5;
  assign state_output_0_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_0_sva,
      or_17_nl);
  assign or_19_nl = or_dcpl_8 | or_dcpl_10;
  assign state_output_1_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_1_sva,
      or_19_nl);
  assign or_22_nl = or_dcpl_13 | or_dcpl_5;
  assign state_output_2_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_2_sva,
      or_22_nl);
  assign or_23_nl = or_dcpl_13 | or_dcpl_10;
  assign state_output_3_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_3_sva,
      or_23_nl);
  assign or_26_nl = or_dcpl_17 | or_dcpl_5;
  assign state_output_4_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_4_sva,
      or_26_nl);
  assign or_27_nl = or_dcpl_17 | or_dcpl_10;
  assign state_output_5_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_5_sva,
      or_27_nl);
  assign or_30_nl = or_dcpl_21 | or_dcpl_5;
  assign state_output_6_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_6_sva,
      or_30_nl);
  assign or_31_nl = or_dcpl_21 | or_dcpl_10;
  assign state_output_7_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_7_sva,
      or_31_nl);
  assign or_34_nl = or_dcpl_8 | or_dcpl_25;
  assign state_output_8_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_8_sva,
      or_34_nl);
  assign or_36_nl = or_dcpl_8 | or_dcpl_27;
  assign state_output_9_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_9_sva,
      or_36_nl);
  assign or_37_nl = or_dcpl_13 | or_dcpl_25;
  assign state_output_10_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_10_sva,
      or_37_nl);
  assign or_38_nl = or_dcpl_13 | or_dcpl_27;
  assign state_output_11_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_11_sva,
      or_38_nl);
  assign or_39_nl = or_dcpl_17 | or_dcpl_25;
  assign state_output_12_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_12_sva,
      or_39_nl);
  assign or_40_nl = or_dcpl_17 | or_dcpl_27;
  assign state_output_13_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_13_sva,
      or_40_nl);
  assign or_41_nl = or_dcpl_21 | or_dcpl_25;
  assign state_output_14_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_14_sva,
      or_41_nl);
  assign or_42_nl = or_dcpl_21 | or_dcpl_27;
  assign state_output_15_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_15_sva,
      or_42_nl);
  assign or_45_nl = or_dcpl_36 | or_dcpl_5;
  assign state_output_16_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_16_sva,
      or_45_nl);
  assign or_46_nl = or_dcpl_36 | or_dcpl_10;
  assign state_output_17_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_17_sva,
      or_46_nl);
  assign or_48_nl = or_dcpl_39 | or_dcpl_5;
  assign state_output_18_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_18_sva,
      or_48_nl);
  assign or_49_nl = or_dcpl_39 | or_dcpl_10;
  assign state_output_19_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_19_sva,
      or_49_nl);
  assign or_51_nl = or_dcpl_42 | or_dcpl_5;
  assign state_output_20_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_20_sva,
      or_51_nl);
  assign or_52_nl = or_dcpl_42 | or_dcpl_10;
  assign state_output_21_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_21_sva,
      or_52_nl);
  assign or_54_nl = or_dcpl_45 | or_dcpl_5;
  assign state_output_22_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_22_sva,
      or_54_nl);
  assign or_55_nl = or_dcpl_45 | or_dcpl_10;
  assign state_output_23_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_23_sva,
      or_55_nl);
  assign or_56_nl = or_dcpl_36 | or_dcpl_25;
  assign state_output_24_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_24_sva,
      or_56_nl);
  assign or_57_nl = or_dcpl_36 | or_dcpl_27;
  assign state_output_25_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_25_sva,
      or_57_nl);
  assign or_58_nl = or_dcpl_39 | or_dcpl_25;
  assign state_output_26_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_26_sva,
      or_58_nl);
  assign or_59_nl = or_dcpl_39 | or_dcpl_27;
  assign state_output_27_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_27_sva,
      or_59_nl);
  assign or_60_nl = or_dcpl_42 | or_dcpl_25;
  assign state_output_28_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_28_sva,
      or_60_nl);
  assign or_61_nl = or_dcpl_42 | or_dcpl_27;
  assign state_output_29_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_29_sva,
      or_61_nl);
  assign or_62_nl = or_dcpl_45 | or_dcpl_25;
  assign state_output_30_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_30_sva,
      or_62_nl);
  assign or_63_nl = or_dcpl_45 | or_dcpl_27;
  assign state_output_31_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_31_sva,
      or_63_nl);
  assign or_66_nl = or_dcpl_57 | or_dcpl_5;
  assign state_output_32_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_32_sva,
      or_66_nl);
  assign or_67_nl = or_dcpl_57 | or_dcpl_10;
  assign state_output_33_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_33_sva,
      or_67_nl);
  assign or_69_nl = or_dcpl_60 | or_dcpl_5;
  assign state_output_34_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_34_sva,
      or_69_nl);
  assign or_70_nl = or_dcpl_60 | or_dcpl_10;
  assign state_output_35_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_35_sva,
      or_70_nl);
  assign or_72_nl = or_dcpl_63 | or_dcpl_5;
  assign state_output_36_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_36_sva,
      or_72_nl);
  assign or_73_nl = or_dcpl_63 | or_dcpl_10;
  assign state_output_37_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_37_sva,
      or_73_nl);
  assign or_75_nl = or_dcpl_66 | or_dcpl_5;
  assign state_output_38_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_38_sva,
      or_75_nl);
  assign or_76_nl = or_dcpl_66 | or_dcpl_10;
  assign state_output_39_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_39_sva,
      or_76_nl);
  assign or_77_nl = or_dcpl_57 | or_dcpl_25;
  assign state_output_40_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_40_sva,
      or_77_nl);
  assign or_78_nl = or_dcpl_57 | or_dcpl_27;
  assign state_output_41_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_41_sva,
      or_78_nl);
  assign or_79_nl = or_dcpl_60 | or_dcpl_25;
  assign state_output_42_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_42_sva,
      or_79_nl);
  assign or_80_nl = or_dcpl_60 | or_dcpl_27;
  assign state_output_43_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_43_sva,
      or_80_nl);
  assign or_81_nl = or_dcpl_63 | or_dcpl_25;
  assign state_output_44_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_44_sva,
      or_81_nl);
  assign or_82_nl = or_dcpl_63 | or_dcpl_27;
  assign state_output_45_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_45_sva,
      or_82_nl);
  assign or_83_nl = or_dcpl_66 | or_dcpl_25;
  assign state_output_46_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_46_sva,
      or_83_nl);
  assign or_84_nl = or_dcpl_66 | or_dcpl_27;
  assign state_output_47_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_47_sva,
      or_84_nl);
  assign or_87_nl = or_dcpl_78 | or_dcpl_5;
  assign state_output_48_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_48_sva,
      or_87_nl);
  assign or_88_nl = or_dcpl_78 | or_dcpl_10;
  assign state_output_49_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_49_sva,
      or_88_nl);
  assign or_90_nl = or_dcpl_81 | or_dcpl_5;
  assign state_output_50_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_50_sva,
      or_90_nl);
  assign or_91_nl = or_dcpl_81 | or_dcpl_10;
  assign state_output_51_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_51_sva,
      or_91_nl);
  assign or_93_nl = or_dcpl_84 | or_dcpl_5;
  assign state_output_52_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_52_sva,
      or_93_nl);
  assign or_94_nl = or_dcpl_84 | or_dcpl_10;
  assign state_output_53_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_53_sva,
      or_94_nl);
  assign or_96_nl = or_dcpl_87 | or_dcpl_5;
  assign state_output_54_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_54_sva,
      or_96_nl);
  assign or_97_nl = or_dcpl_87 | or_dcpl_10;
  assign state_output_55_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_55_sva,
      or_97_nl);
  assign or_98_nl = or_dcpl_78 | or_dcpl_25;
  assign state_output_56_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_56_sva,
      or_98_nl);
  assign or_99_nl = or_dcpl_78 | or_dcpl_27;
  assign state_output_57_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_57_sva,
      or_99_nl);
  assign or_100_nl = or_dcpl_81 | or_dcpl_25;
  assign state_output_58_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_58_sva,
      or_100_nl);
  assign or_101_nl = or_dcpl_81 | or_dcpl_27;
  assign state_output_59_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_59_sva,
      or_101_nl);
  assign or_102_nl = or_dcpl_84 | or_dcpl_25;
  assign state_output_60_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_60_sva,
      or_102_nl);
  assign or_103_nl = or_dcpl_84 | or_dcpl_27;
  assign state_output_61_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_61_sva,
      or_103_nl);
  assign or_104_nl = or_dcpl_87 | or_dcpl_25;
  assign state_output_62_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_62_sva,
      or_104_nl);
  assign or_105_nl = or_dcpl_87 | or_dcpl_27;
  assign state_output_63_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_63_sva,
      or_105_nl);
  assign or_108_nl = or_dcpl_8 | or_dcpl_99;
  assign state_output_64_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_64_sva,
      or_108_nl);
  assign or_110_nl = or_dcpl_8 | or_dcpl_101;
  assign state_output_65_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_65_sva,
      or_110_nl);
  assign or_111_nl = or_dcpl_13 | or_dcpl_99;
  assign state_output_66_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_66_sva,
      or_111_nl);
  assign or_112_nl = or_dcpl_13 | or_dcpl_101;
  assign state_output_67_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_67_sva,
      or_112_nl);
  assign or_113_nl = or_dcpl_17 | or_dcpl_99;
  assign state_output_68_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_68_sva,
      or_113_nl);
  assign or_114_nl = or_dcpl_17 | or_dcpl_101;
  assign state_output_69_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_69_sva,
      or_114_nl);
  assign or_115_nl = or_dcpl_21 | or_dcpl_99;
  assign state_output_70_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_70_sva,
      or_115_nl);
  assign or_116_nl = or_dcpl_21 | or_dcpl_101;
  assign state_output_71_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_71_sva,
      or_116_nl);
  assign or_119_nl = or_dcpl_8 | or_dcpl_110;
  assign state_output_72_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_72_sva,
      or_119_nl);
  assign or_121_nl = or_dcpl_8 | or_dcpl_112;
  assign state_output_73_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_73_sva,
      or_121_nl);
  assign or_122_nl = or_dcpl_13 | or_dcpl_110;
  assign state_output_74_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_74_sva,
      or_122_nl);
  assign or_123_nl = or_dcpl_13 | or_dcpl_112;
  assign state_output_75_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_75_sva,
      or_123_nl);
  assign or_124_nl = or_dcpl_17 | or_dcpl_110;
  assign state_output_76_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_76_sva,
      or_124_nl);
  assign or_125_nl = or_dcpl_17 | or_dcpl_112;
  assign state_output_77_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_77_sva,
      or_125_nl);
  assign or_126_nl = or_dcpl_21 | or_dcpl_110;
  assign state_output_78_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_78_sva,
      or_126_nl);
  assign or_127_nl = or_dcpl_21 | or_dcpl_112;
  assign state_output_79_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_79_sva,
      or_127_nl);
  assign or_128_nl = or_dcpl_36 | or_dcpl_99;
  assign state_output_80_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_80_sva,
      or_128_nl);
  assign or_129_nl = or_dcpl_36 | or_dcpl_101;
  assign state_output_81_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_81_sva,
      or_129_nl);
  assign or_130_nl = or_dcpl_39 | or_dcpl_99;
  assign state_output_82_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_82_sva,
      or_130_nl);
  assign or_131_nl = or_dcpl_39 | or_dcpl_101;
  assign state_output_83_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_83_sva,
      or_131_nl);
  assign or_132_nl = or_dcpl_42 | or_dcpl_99;
  assign state_output_84_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_84_sva,
      or_132_nl);
  assign or_133_nl = or_dcpl_42 | or_dcpl_101;
  assign state_output_85_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_85_sva,
      or_133_nl);
  assign or_134_nl = or_dcpl_45 | or_dcpl_99;
  assign state_output_86_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_86_sva,
      or_134_nl);
  assign or_135_nl = or_dcpl_45 | or_dcpl_101;
  assign state_output_87_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_87_sva,
      or_135_nl);
  assign or_136_nl = or_dcpl_36 | or_dcpl_110;
  assign state_output_88_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_88_sva,
      or_136_nl);
  assign or_137_nl = or_dcpl_36 | or_dcpl_112;
  assign state_output_89_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_89_sva,
      or_137_nl);
  assign or_138_nl = or_dcpl_39 | or_dcpl_110;
  assign state_output_90_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_90_sva,
      or_138_nl);
  assign or_139_nl = or_dcpl_39 | or_dcpl_112;
  assign state_output_91_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_91_sva,
      or_139_nl);
  assign or_140_nl = or_dcpl_42 | or_dcpl_110;
  assign state_output_92_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_92_sva,
      or_140_nl);
  assign or_141_nl = or_dcpl_42 | or_dcpl_112;
  assign state_output_93_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_93_sva,
      or_141_nl);
  assign or_142_nl = or_dcpl_45 | or_dcpl_110;
  assign state_output_94_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_94_sva,
      or_142_nl);
  assign or_143_nl = or_dcpl_45 | or_dcpl_112;
  assign state_output_95_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_95_sva,
      or_143_nl);
  assign or_144_nl = or_dcpl_57 | or_dcpl_99;
  assign state_output_96_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_96_sva,
      or_144_nl);
  assign or_145_nl = or_dcpl_57 | or_dcpl_101;
  assign state_output_97_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_97_sva,
      or_145_nl);
  assign or_146_nl = or_dcpl_60 | or_dcpl_99;
  assign state_output_98_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_98_sva,
      or_146_nl);
  assign or_147_nl = or_dcpl_60 | or_dcpl_101;
  assign state_output_99_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_99_sva,
      or_147_nl);
  assign or_148_nl = or_dcpl_63 | or_dcpl_99;
  assign state_output_100_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_100_sva,
      or_148_nl);
  assign or_149_nl = or_dcpl_63 | or_dcpl_101;
  assign state_output_101_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_101_sva,
      or_149_nl);
  assign or_150_nl = or_dcpl_66 | or_dcpl_99;
  assign state_output_102_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_102_sva,
      or_150_nl);
  assign or_151_nl = or_dcpl_66 | or_dcpl_101;
  assign state_output_103_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_103_sva,
      or_151_nl);
  assign or_152_nl = or_dcpl_57 | or_dcpl_110;
  assign state_output_104_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_104_sva,
      or_152_nl);
  assign or_153_nl = or_dcpl_57 | or_dcpl_112;
  assign state_output_105_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_105_sva,
      or_153_nl);
  assign or_154_nl = or_dcpl_60 | or_dcpl_110;
  assign state_output_106_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_106_sva,
      or_154_nl);
  assign or_155_nl = or_dcpl_60 | or_dcpl_112;
  assign state_output_107_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_107_sva,
      or_155_nl);
  assign or_156_nl = or_dcpl_63 | or_dcpl_110;
  assign state_output_108_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_108_sva,
      or_156_nl);
  assign or_157_nl = or_dcpl_63 | or_dcpl_112;
  assign state_output_109_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_109_sva,
      or_157_nl);
  assign or_158_nl = or_dcpl_66 | or_dcpl_110;
  assign state_output_110_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_110_sva,
      or_158_nl);
  assign or_159_nl = or_dcpl_66 | or_dcpl_112;
  assign state_output_111_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_111_sva,
      or_159_nl);
  assign or_160_nl = or_dcpl_78 | or_dcpl_99;
  assign state_output_112_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_112_sva,
      or_160_nl);
  assign or_161_nl = or_dcpl_78 | or_dcpl_101;
  assign state_output_113_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_113_sva,
      or_161_nl);
  assign or_162_nl = or_dcpl_81 | or_dcpl_99;
  assign state_output_114_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_114_sva,
      or_162_nl);
  assign or_163_nl = or_dcpl_81 | or_dcpl_101;
  assign state_output_115_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_115_sva,
      or_163_nl);
  assign or_164_nl = or_dcpl_84 | or_dcpl_99;
  assign state_output_116_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_116_sva,
      or_164_nl);
  assign or_165_nl = or_dcpl_84 | or_dcpl_101;
  assign state_output_117_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_117_sva,
      or_165_nl);
  assign or_166_nl = or_dcpl_87 | or_dcpl_99;
  assign state_output_118_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_118_sva,
      or_166_nl);
  assign or_167_nl = or_dcpl_87 | or_dcpl_101;
  assign state_output_119_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_119_sva,
      or_167_nl);
  assign or_168_nl = or_dcpl_78 | or_dcpl_110;
  assign state_output_120_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_120_sva,
      or_168_nl);
  assign or_169_nl = or_dcpl_78 | or_dcpl_112;
  assign state_output_121_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_121_sva,
      or_169_nl);
  assign or_170_nl = or_dcpl_81 | or_dcpl_110;
  assign state_output_122_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_122_sva,
      or_170_nl);
  assign or_171_nl = or_dcpl_81 | or_dcpl_112;
  assign state_output_123_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_123_sva,
      or_171_nl);
  assign or_172_nl = or_dcpl_84 | or_dcpl_110;
  assign state_output_124_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_124_sva,
      or_172_nl);
  assign or_173_nl = or_dcpl_84 | or_dcpl_112;
  assign state_output_125_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_125_sva,
      or_173_nl);
  assign or_174_nl = or_dcpl_87 | or_dcpl_110;
  assign state_output_126_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_126_sva,
      or_174_nl);
  assign or_175_nl = or_dcpl_87 | or_dcpl_112;
  assign state_output_127_sva_1_mx0 = MUX_v_16_2_2(acc_out_rsci_idat, state_output_127_sva,
      or_175_nl);
  assign aqed_in_if_mux_7_nl = MUX_s_1_2_2(state_orig_idx_sva, (~ original_rsci_idat),
      aqed_in_if_issue_orig_land_lpi_1_dfm_1);
  assign state_orig_idx_sva_dfm_1_mx0 = MUX_s_1_2_2(state_orig_idx_sva, (aqed_in_if_mux_7_nl),
      bmc_v_rsci_idat);
  assign state_dup_in_sva_dfm_1_mx0 = MUX_v_16_2_2(state_in_count_sva, state_dup_in_sva,
      state_dup_issued_sva);
  assign aqed_in_if_mux_8_nl = MUX_s_1_2_2(state_dup_idx_sva, (~ duplicate_rsci_idat),
      aqed_in_if_issue_dup_land_1_lpi_1_dfm_2);
  assign state_dup_idx_sva_dfm_1_mx0 = MUX_s_1_2_2(state_dup_idx_sva, (aqed_in_if_mux_8_nl),
      bmc_v_rsci_idat);
  assign and_9_cse = original_rsci_idat & bmc_v_rsci_idat;
  assign nl_aqed_out_if_aelse_2_acc_nl = ({1'b1 , state_out_count_sva}) + conv_u2u_16_17(~
      state_dup_in_sva_dfm_1_mx0) + 17'b00000000000000001;
  assign aqed_out_if_aelse_2_acc_nl = nl_aqed_out_if_aelse_2_acc_nl[16:0];
  assign aqed_out_if_aelse_2_acc_itm_16 = readslicef_17_1_16((aqed_out_if_aelse_2_acc_nl));
  assign aqed_in_if_issue_dup_land_1_lpi_1_dfm_2 = (aqed_in_if_issue_orig_land_lpi_1_dfm_1
      | (aqed_in_if_issue_dup_aif_1_aif_equal_tmp & state_orig_issued_sva)) & (~
      state_dup_issued_sva) & duplicate_rsci_idat;
  assign aqed_in_if_issue_orig_land_lpi_1_dfm_1 = (~ state_orig_issued_sva) & original_rsci_idat;
  assign aqed_in_if_issue_dup_aif_1_aif_equal_tmp = bmc_in_rsci_idat == state_dup_in_sva;
  assign aqed_in_if_aqed_in_if_or_2_nl = state_orig_issued_sva | aqed_in_if_issue_orig_land_lpi_1_dfm_1;
  assign state_orig_issued_sva_mx0 = MUX_s_1_2_2(state_orig_issued_sva, (aqed_in_if_aqed_in_if_or_2_nl),
      bmc_v_rsci_idat);
  assign aqed_in_if_aqed_in_if_or_3_nl = state_dup_issued_sva | aqed_in_if_issue_dup_land_1_lpi_1_dfm_2;
  assign state_dup_issued_sva_mx0 = MUX_s_1_2_2(state_dup_issued_sva, (aqed_in_if_aqed_in_if_or_3_nl),
      bmc_v_rsci_idat);
  assign aqed_out_if_aqed_out_if_and_1_tmp = acc_out_rdy_rsci_idat & acc_out_v_rsci_idat;
  assign and_dcpl = ~((~((~ mux_6_cse) | aqed_out_if_aelse_2_acc_itm_16 | (~ aqed_out_if_aqed_out_if_and_1_tmp)))
      | state_qed_done_sva);
  assign or_dcpl_4 = (state_out_count_sva[3]) | (state_out_count_sva[6]);
  assign or_dcpl_5 = or_dcpl_4 | (state_out_count_sva[0]);
  assign or_dcpl_6 = (state_out_count_sva[2:1]!=2'b00);
  assign or_dcpl_7 = (state_out_count_sva[5:4]!=2'b00);
  assign or_dcpl_8 = or_dcpl_7 | or_dcpl_6;
  assign or_dcpl_10 = or_dcpl_4 | (~ (state_out_count_sva[0]));
  assign or_dcpl_12 = (state_out_count_sva[2:1]!=2'b01);
  assign or_dcpl_13 = or_dcpl_7 | or_dcpl_12;
  assign or_dcpl_16 = (state_out_count_sva[2:1]!=2'b10);
  assign or_dcpl_17 = or_dcpl_7 | or_dcpl_16;
  assign or_dcpl_20 = ~((state_out_count_sva[2:1]==2'b11));
  assign or_dcpl_21 = or_dcpl_7 | or_dcpl_20;
  assign or_dcpl_24 = (~ (state_out_count_sva[3])) | (state_out_count_sva[6]);
  assign or_dcpl_25 = or_dcpl_24 | (state_out_count_sva[0]);
  assign or_dcpl_27 = or_dcpl_24 | (~ (state_out_count_sva[0]));
  assign or_dcpl_35 = (state_out_count_sva[5:4]!=2'b01);
  assign or_dcpl_36 = or_dcpl_35 | or_dcpl_6;
  assign or_dcpl_39 = or_dcpl_35 | or_dcpl_12;
  assign or_dcpl_42 = or_dcpl_35 | or_dcpl_16;
  assign or_dcpl_45 = or_dcpl_35 | or_dcpl_20;
  assign or_dcpl_56 = (state_out_count_sva[5:4]!=2'b10);
  assign or_dcpl_57 = or_dcpl_56 | or_dcpl_6;
  assign or_dcpl_60 = or_dcpl_56 | or_dcpl_12;
  assign or_dcpl_63 = or_dcpl_56 | or_dcpl_16;
  assign or_dcpl_66 = or_dcpl_56 | or_dcpl_20;
  assign or_dcpl_77 = ~((state_out_count_sva[5:4]==2'b11));
  assign or_dcpl_78 = or_dcpl_77 | or_dcpl_6;
  assign or_dcpl_81 = or_dcpl_77 | or_dcpl_12;
  assign or_dcpl_84 = or_dcpl_77 | or_dcpl_16;
  assign or_dcpl_87 = or_dcpl_77 | or_dcpl_20;
  assign or_dcpl_98 = (state_out_count_sva[3]) | (~ (state_out_count_sva[6]));
  assign or_dcpl_99 = or_dcpl_98 | (state_out_count_sva[0]);
  assign or_dcpl_101 = or_dcpl_98 | (~ (state_out_count_sva[0]));
  assign or_dcpl_109 = ~((state_out_count_sva[3]) & (state_out_count_sva[6]));
  assign or_dcpl_110 = or_dcpl_109 | (state_out_count_sva[0]);
  assign or_dcpl_112 = or_dcpl_109 | (~ (state_out_count_sva[0]));
  assign or_dcpl_168 = ~((state_out_count_sva[0]) & aqed_out_if_aqed_out_if_and_1_tmp);
  assign or_dcpl_169 = or_dcpl_24 | or_dcpl_168;
  assign or_dcpl_171 = (state_out_count_sva[0]) | (~ aqed_out_if_aqed_out_if_and_1_tmp);
  assign or_dcpl_172 = or_dcpl_98 | or_dcpl_171;
  assign or_dcpl_174 = or_dcpl_24 | or_dcpl_171;
  assign or_dcpl_176 = or_dcpl_98 | or_dcpl_168;
  assign or_dcpl_190 = or_dcpl_4 | or_dcpl_168;
  assign or_dcpl_192 = or_dcpl_109 | or_dcpl_171;
  assign or_dcpl_194 = or_dcpl_4 | or_dcpl_171;
  assign or_dcpl_196 = or_dcpl_109 | or_dcpl_168;
  assign and_dcpl_23 = bmc_v_rsci_idat & clk_en;
  always @(posedge clk) begin
    if ( reset ) begin
      state_out_count_sva <= 16'b0000000000000000;
      state_qed_done_sva <= 1'b0;
      reg_state_orig_done_cse <= 1'b0;
    end
    else if ( state_out_count_and_cse ) begin
      state_out_count_sva <= nl_state_out_count_sva[15:0];
      state_qed_done_sva <= state_qed_done_sva | ((~ aqed_out_if_aelse_2_acc_itm_16)
          & state_dup_issued_sva_mx0 & state_orig_issued_sva_mx0);
      reg_state_orig_done_cse <= (~ (readslicef_17_1_16((aqed_out_if_aelse_acc_nl))))
          & state_orig_issued_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_63_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_169)) ) begin
      state_output_63_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_64_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_172)) ) begin
      state_output_64_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_62_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_174)) ) begin
      state_output_62_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_65_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_176)) ) begin
      state_output_65_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_61_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_169)) ) begin
      state_output_61_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_66_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_172)) ) begin
      state_output_66_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_60_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_174)) ) begin
      state_output_60_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_67_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_176)) ) begin
      state_output_67_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_59_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_169)) ) begin
      state_output_59_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_68_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_172)) ) begin
      state_output_68_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_58_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_174)) ) begin
      state_output_58_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_69_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_176)) ) begin
      state_output_69_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_57_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_169)) ) begin
      state_output_57_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_70_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_172)) ) begin
      state_output_70_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_56_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_174)) ) begin
      state_output_56_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_71_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_176)) ) begin
      state_output_71_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_55_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_190)) ) begin
      state_output_55_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_72_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_192)) ) begin
      state_output_72_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_54_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_194)) ) begin
      state_output_54_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_73_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_196)) ) begin
      state_output_73_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_53_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_190)) ) begin
      state_output_53_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_74_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_192)) ) begin
      state_output_74_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_52_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_194)) ) begin
      state_output_52_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_75_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_196)) ) begin
      state_output_75_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_51_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_190)) ) begin
      state_output_51_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_76_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_192)) ) begin
      state_output_76_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_50_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_194)) ) begin
      state_output_50_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_77_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_196)) ) begin
      state_output_77_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_49_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_190)) ) begin
      state_output_49_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_78_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_192)) ) begin
      state_output_78_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_48_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_194)) ) begin
      state_output_48_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_79_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_196)) ) begin
      state_output_79_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_47_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_169)) ) begin
      state_output_47_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_80_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_172)) ) begin
      state_output_80_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_46_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_174)) ) begin
      state_output_46_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_81_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_176)) ) begin
      state_output_81_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_45_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_169)) ) begin
      state_output_45_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_82_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_172)) ) begin
      state_output_82_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_44_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_174)) ) begin
      state_output_44_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_83_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_176)) ) begin
      state_output_83_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_43_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_169)) ) begin
      state_output_43_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_84_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_172)) ) begin
      state_output_84_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_42_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_174)) ) begin
      state_output_42_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_85_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_176)) ) begin
      state_output_85_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_41_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_169)) ) begin
      state_output_41_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_86_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_172)) ) begin
      state_output_86_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_40_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_174)) ) begin
      state_output_40_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_87_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_176)) ) begin
      state_output_87_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_39_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_190)) ) begin
      state_output_39_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_88_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_192)) ) begin
      state_output_88_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_38_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_194)) ) begin
      state_output_38_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_89_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_196)) ) begin
      state_output_89_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_37_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_190)) ) begin
      state_output_37_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_90_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_192)) ) begin
      state_output_90_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_36_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_194)) ) begin
      state_output_36_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_91_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_196)) ) begin
      state_output_91_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_35_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_190)) ) begin
      state_output_35_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_92_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_192)) ) begin
      state_output_92_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_34_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_194)) ) begin
      state_output_34_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_93_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_196)) ) begin
      state_output_93_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_33_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_190)) ) begin
      state_output_33_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_94_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_192)) ) begin
      state_output_94_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_32_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_194)) ) begin
      state_output_32_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_95_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_196)) ) begin
      state_output_95_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_31_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_169)) ) begin
      state_output_31_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_96_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_172)) ) begin
      state_output_96_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_30_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_174)) ) begin
      state_output_30_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_97_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_176)) ) begin
      state_output_97_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_29_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_169)) ) begin
      state_output_29_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_98_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_172)) ) begin
      state_output_98_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_28_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_174)) ) begin
      state_output_28_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_99_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_176)) ) begin
      state_output_99_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_27_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_169)) ) begin
      state_output_27_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_100_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_172)) ) begin
      state_output_100_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_26_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_174)) ) begin
      state_output_26_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_101_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_176)) ) begin
      state_output_101_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_25_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_169)) ) begin
      state_output_25_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_102_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_172)) ) begin
      state_output_102_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_24_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_174)) ) begin
      state_output_24_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_103_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_176)) ) begin
      state_output_103_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_23_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_190)) ) begin
      state_output_23_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_104_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_192)) ) begin
      state_output_104_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_22_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_45 | or_dcpl_194)) ) begin
      state_output_22_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_105_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_57 | or_dcpl_196)) ) begin
      state_output_105_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_21_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_190)) ) begin
      state_output_21_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_106_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_192)) ) begin
      state_output_106_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_20_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_42 | or_dcpl_194)) ) begin
      state_output_20_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_107_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_60 | or_dcpl_196)) ) begin
      state_output_107_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_19_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_190)) ) begin
      state_output_19_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_108_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_192)) ) begin
      state_output_108_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_18_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_39 | or_dcpl_194)) ) begin
      state_output_18_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_109_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_63 | or_dcpl_196)) ) begin
      state_output_109_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_17_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_190)) ) begin
      state_output_17_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_110_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_192)) ) begin
      state_output_110_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_16_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_36 | or_dcpl_194)) ) begin
      state_output_16_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_111_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_66 | or_dcpl_196)) ) begin
      state_output_111_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_15_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_169)) ) begin
      state_output_15_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_112_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_172)) ) begin
      state_output_112_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_14_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_174)) ) begin
      state_output_14_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_113_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_176)) ) begin
      state_output_113_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_13_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_169)) ) begin
      state_output_13_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_114_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_172)) ) begin
      state_output_114_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_12_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_174)) ) begin
      state_output_12_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_115_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_176)) ) begin
      state_output_115_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_11_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_169)) ) begin
      state_output_11_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_116_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_172)) ) begin
      state_output_116_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_10_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_174)) ) begin
      state_output_10_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_117_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_176)) ) begin
      state_output_117_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_9_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_169)) ) begin
      state_output_9_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_118_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_172)) ) begin
      state_output_118_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_8_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_174)) ) begin
      state_output_8_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_119_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_176)) ) begin
      state_output_119_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_7_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_190)) ) begin
      state_output_7_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_120_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_192)) ) begin
      state_output_120_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_6_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_21 | or_dcpl_194)) ) begin
      state_output_6_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_121_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_78 | or_dcpl_196)) ) begin
      state_output_121_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_5_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_190)) ) begin
      state_output_5_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_122_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_192)) ) begin
      state_output_122_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_4_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_17 | or_dcpl_194)) ) begin
      state_output_4_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_123_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_81 | or_dcpl_196)) ) begin
      state_output_123_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_3_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_190)) ) begin
      state_output_3_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_124_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_192)) ) begin
      state_output_124_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_2_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_13 | or_dcpl_194)) ) begin
      state_output_2_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_125_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_84 | or_dcpl_196)) ) begin
      state_output_125_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_1_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_190)) ) begin
      state_output_1_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_126_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_192)) ) begin
      state_output_126_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_0_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_8 | or_dcpl_194)) ) begin
      state_output_0_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_output_127_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & and_dcpl & (~(or_dcpl_87 | or_dcpl_196)) ) begin
      state_output_127_sva <= acc_out_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      reg_state_qed_check_cse <= 1'b0;
    end
    else if ( clk_en & (~((~ mux_6_cse) | aqed_out_if_aelse_2_acc_itm_16 | (~ aqed_out_if_aqed_out_if_and_1_tmp)
        | state_qed_done_sva)) ) begin
      reg_state_qed_check_cse <= (aqed_out_if_if_mux_nl) == (aqed_out_if_if_mux_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_dup_idx_sva <= 1'b0;
    end
    else if ( (mux_nl) & ((~(acc_out_v_rsci_idat & acc_out_rdy_rsci_idat)) | aqed_out_if_aelse_2_acc_itm_16)
        & clk_en & (~ state_qed_done_sva) & duplicate_rsci_idat & bmc_v_rsci_idat
        & (~ state_dup_issued_sva) ) begin
      state_dup_idx_sva <= state_dup_idx_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_idx_sva <= 1'b0;
    end
    else if ( ((~((duplicate_rsci_idat | state_dup_issued_sva) & acc_out_v_rsci_idat))
        | (~ acc_out_rdy_rsci_idat) | aqed_out_if_aelse_2_acc_itm_16) & clk_en &
        (~ state_qed_done_sva) & bmc_v_rsci_idat & original_rsci_idat & (~ state_orig_issued_sva)
        ) begin
      state_orig_idx_sva <= state_orig_idx_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_dup_in_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & (and_9_cse | state_orig_issued_sva | state_dup_issued_sva)
        & (((aqed_in_if_issue_dup_aif_1_aif_equal_tmp | (~ state_orig_issued_sva))
        & bmc_v_rsci_idat & duplicate_rsci_idat & (~ state_dup_issued_sva)) | nor_10_rgt)
        ) begin
      state_dup_in_sva <= MUX_v_16_2_2(state_in_count_sva, bmc_in_rsci_idat, nor_10_rgt);
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_in_count_sva <= 16'b0000000000000000;
    end
    else if ( clk_en & (~ mux_6_cse) & bmc_v_rsci_idat ) begin
      state_in_count_sva <= nl_state_in_count_sva[15:0];
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_in_sva <= 16'b0000000000000000;
    end
    else if ( and_9_cse & (~ state_orig_issued_sva) & clk_en ) begin
      state_orig_in_sva <= state_orig_in_sva_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      state_orig_issued_sva <= 1'b0;
      state_dup_issued_sva <= 1'b0;
    end
    else if ( and_dcpl_23 ) begin
      state_orig_issued_sva <= state_orig_issued_sva_mx0;
      state_dup_issued_sva <= state_dup_issued_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( reset ) begin
      return_aqed_out_v_rsci_idat <= 1'b0;
      return_aqed_out_rsci_idat <= 16'b0000000000000000;
    end
    else if ( clk_en ) begin
      return_aqed_out_v_rsci_idat <= bmc_v_rsci_idat;
      return_aqed_out_rsci_idat <= bmc_in_rsci_idat;
    end
  end
  assign nl_state_out_count_sva  = state_out_count_sva + 16'b0000000000000001;
  assign nl_aqed_out_if_aelse_acc_nl = ({1'b1 , state_out_count_sva}) + conv_u2u_16_17(~
      state_orig_in_sva_dfm_1_mx0) + 17'b00000000000000001;
  assign aqed_out_if_aelse_acc_nl = nl_aqed_out_if_aelse_acc_nl[16:0];
  assign nl_operator_ac_int_16_false_1_false_2_acc_nl = (state_orig_in_sva_dfm_1_mx0[6:0])
      + conv_u2u_1_7(state_orig_idx_sva_dfm_1_mx0);
  assign operator_ac_int_16_false_1_false_2_acc_nl = nl_operator_ac_int_16_false_1_false_2_acc_nl[6:0];
  assign aqed_out_if_if_mux_nl = MUX_v_16_128_2(state_output_0_sva_1_mx0, state_output_1_sva_1_mx0,
      state_output_2_sva_1_mx0, state_output_3_sva_1_mx0, state_output_4_sva_1_mx0,
      state_output_5_sva_1_mx0, state_output_6_sva_1_mx0, state_output_7_sva_1_mx0,
      state_output_8_sva_1_mx0, state_output_9_sva_1_mx0, state_output_10_sva_1_mx0,
      state_output_11_sva_1_mx0, state_output_12_sva_1_mx0, state_output_13_sva_1_mx0,
      state_output_14_sva_1_mx0, state_output_15_sva_1_mx0, state_output_16_sva_1_mx0,
      state_output_17_sva_1_mx0, state_output_18_sva_1_mx0, state_output_19_sva_1_mx0,
      state_output_20_sva_1_mx0, state_output_21_sva_1_mx0, state_output_22_sva_1_mx0,
      state_output_23_sva_1_mx0, state_output_24_sva_1_mx0, state_output_25_sva_1_mx0,
      state_output_26_sva_1_mx0, state_output_27_sva_1_mx0, state_output_28_sva_1_mx0,
      state_output_29_sva_1_mx0, state_output_30_sva_1_mx0, state_output_31_sva_1_mx0,
      state_output_32_sva_1_mx0, state_output_33_sva_1_mx0, state_output_34_sva_1_mx0,
      state_output_35_sva_1_mx0, state_output_36_sva_1_mx0, state_output_37_sva_1_mx0,
      state_output_38_sva_1_mx0, state_output_39_sva_1_mx0, state_output_40_sva_1_mx0,
      state_output_41_sva_1_mx0, state_output_42_sva_1_mx0, state_output_43_sva_1_mx0,
      state_output_44_sva_1_mx0, state_output_45_sva_1_mx0, state_output_46_sva_1_mx0,
      state_output_47_sva_1_mx0, state_output_48_sva_1_mx0, state_output_49_sva_1_mx0,
      state_output_50_sva_1_mx0, state_output_51_sva_1_mx0, state_output_52_sva_1_mx0,
      state_output_53_sva_1_mx0, state_output_54_sva_1_mx0, state_output_55_sva_1_mx0,
      state_output_56_sva_1_mx0, state_output_57_sva_1_mx0, state_output_58_sva_1_mx0,
      state_output_59_sva_1_mx0, state_output_60_sva_1_mx0, state_output_61_sva_1_mx0,
      state_output_62_sva_1_mx0, state_output_63_sva_1_mx0, state_output_64_sva_1_mx0,
      state_output_65_sva_1_mx0, state_output_66_sva_1_mx0, state_output_67_sva_1_mx0,
      state_output_68_sva_1_mx0, state_output_69_sva_1_mx0, state_output_70_sva_1_mx0,
      state_output_71_sva_1_mx0, state_output_72_sva_1_mx0, state_output_73_sva_1_mx0,
      state_output_74_sva_1_mx0, state_output_75_sva_1_mx0, state_output_76_sva_1_mx0,
      state_output_77_sva_1_mx0, state_output_78_sva_1_mx0, state_output_79_sva_1_mx0,
      state_output_80_sva_1_mx0, state_output_81_sva_1_mx0, state_output_82_sva_1_mx0,
      state_output_83_sva_1_mx0, state_output_84_sva_1_mx0, state_output_85_sva_1_mx0,
      state_output_86_sva_1_mx0, state_output_87_sva_1_mx0, state_output_88_sva_1_mx0,
      state_output_89_sva_1_mx0, state_output_90_sva_1_mx0, state_output_91_sva_1_mx0,
      state_output_92_sva_1_mx0, state_output_93_sva_1_mx0, state_output_94_sva_1_mx0,
      state_output_95_sva_1_mx0, state_output_96_sva_1_mx0, state_output_97_sva_1_mx0,
      state_output_98_sva_1_mx0, state_output_99_sva_1_mx0, state_output_100_sva_1_mx0,
      state_output_101_sva_1_mx0, state_output_102_sva_1_mx0, state_output_103_sva_1_mx0,
      state_output_104_sva_1_mx0, state_output_105_sva_1_mx0, state_output_106_sva_1_mx0,
      state_output_107_sva_1_mx0, state_output_108_sva_1_mx0, state_output_109_sva_1_mx0,
      state_output_110_sva_1_mx0, state_output_111_sva_1_mx0, state_output_112_sva_1_mx0,
      state_output_113_sva_1_mx0, state_output_114_sva_1_mx0, state_output_115_sva_1_mx0,
      state_output_116_sva_1_mx0, state_output_117_sva_1_mx0, state_output_118_sva_1_mx0,
      state_output_119_sva_1_mx0, state_output_120_sva_1_mx0, state_output_121_sva_1_mx0,
      state_output_122_sva_1_mx0, state_output_123_sva_1_mx0, state_output_124_sva_1_mx0,
      state_output_125_sva_1_mx0, state_output_126_sva_1_mx0, state_output_127_sva_1_mx0,
      operator_ac_int_16_false_1_false_2_acc_nl);
  assign nl_operator_ac_int_16_false_1_false_3_acc_nl = (state_dup_in_sva_dfm_1_mx0[6:0])
      + conv_u2u_1_7(state_dup_idx_sva_dfm_1_mx0);
  assign operator_ac_int_16_false_1_false_3_acc_nl = nl_operator_ac_int_16_false_1_false_3_acc_nl[6:0];
  assign aqed_out_if_if_mux_3_nl = MUX_v_16_128_2(state_output_0_sva_1_mx0, state_output_1_sva_1_mx0,
      state_output_2_sva_1_mx0, state_output_3_sva_1_mx0, state_output_4_sva_1_mx0,
      state_output_5_sva_1_mx0, state_output_6_sva_1_mx0, state_output_7_sva_1_mx0,
      state_output_8_sva_1_mx0, state_output_9_sva_1_mx0, state_output_10_sva_1_mx0,
      state_output_11_sva_1_mx0, state_output_12_sva_1_mx0, state_output_13_sva_1_mx0,
      state_output_14_sva_1_mx0, state_output_15_sva_1_mx0, state_output_16_sva_1_mx0,
      state_output_17_sva_1_mx0, state_output_18_sva_1_mx0, state_output_19_sva_1_mx0,
      state_output_20_sva_1_mx0, state_output_21_sva_1_mx0, state_output_22_sva_1_mx0,
      state_output_23_sva_1_mx0, state_output_24_sva_1_mx0, state_output_25_sva_1_mx0,
      state_output_26_sva_1_mx0, state_output_27_sva_1_mx0, state_output_28_sva_1_mx0,
      state_output_29_sva_1_mx0, state_output_30_sva_1_mx0, state_output_31_sva_1_mx0,
      state_output_32_sva_1_mx0, state_output_33_sva_1_mx0, state_output_34_sva_1_mx0,
      state_output_35_sva_1_mx0, state_output_36_sva_1_mx0, state_output_37_sva_1_mx0,
      state_output_38_sva_1_mx0, state_output_39_sva_1_mx0, state_output_40_sva_1_mx0,
      state_output_41_sva_1_mx0, state_output_42_sva_1_mx0, state_output_43_sva_1_mx0,
      state_output_44_sva_1_mx0, state_output_45_sva_1_mx0, state_output_46_sva_1_mx0,
      state_output_47_sva_1_mx0, state_output_48_sva_1_mx0, state_output_49_sva_1_mx0,
      state_output_50_sva_1_mx0, state_output_51_sva_1_mx0, state_output_52_sva_1_mx0,
      state_output_53_sva_1_mx0, state_output_54_sva_1_mx0, state_output_55_sva_1_mx0,
      state_output_56_sva_1_mx0, state_output_57_sva_1_mx0, state_output_58_sva_1_mx0,
      state_output_59_sva_1_mx0, state_output_60_sva_1_mx0, state_output_61_sva_1_mx0,
      state_output_62_sva_1_mx0, state_output_63_sva_1_mx0, state_output_64_sva_1_mx0,
      state_output_65_sva_1_mx0, state_output_66_sva_1_mx0, state_output_67_sva_1_mx0,
      state_output_68_sva_1_mx0, state_output_69_sva_1_mx0, state_output_70_sva_1_mx0,
      state_output_71_sva_1_mx0, state_output_72_sva_1_mx0, state_output_73_sva_1_mx0,
      state_output_74_sva_1_mx0, state_output_75_sva_1_mx0, state_output_76_sva_1_mx0,
      state_output_77_sva_1_mx0, state_output_78_sva_1_mx0, state_output_79_sva_1_mx0,
      state_output_80_sva_1_mx0, state_output_81_sva_1_mx0, state_output_82_sva_1_mx0,
      state_output_83_sva_1_mx0, state_output_84_sva_1_mx0, state_output_85_sva_1_mx0,
      state_output_86_sva_1_mx0, state_output_87_sva_1_mx0, state_output_88_sva_1_mx0,
      state_output_89_sva_1_mx0, state_output_90_sva_1_mx0, state_output_91_sva_1_mx0,
      state_output_92_sva_1_mx0, state_output_93_sva_1_mx0, state_output_94_sva_1_mx0,
      state_output_95_sva_1_mx0, state_output_96_sva_1_mx0, state_output_97_sva_1_mx0,
      state_output_98_sva_1_mx0, state_output_99_sva_1_mx0, state_output_100_sva_1_mx0,
      state_output_101_sva_1_mx0, state_output_102_sva_1_mx0, state_output_103_sva_1_mx0,
      state_output_104_sva_1_mx0, state_output_105_sva_1_mx0, state_output_106_sva_1_mx0,
      state_output_107_sva_1_mx0, state_output_108_sva_1_mx0, state_output_109_sva_1_mx0,
      state_output_110_sva_1_mx0, state_output_111_sva_1_mx0, state_output_112_sva_1_mx0,
      state_output_113_sva_1_mx0, state_output_114_sva_1_mx0, state_output_115_sva_1_mx0,
      state_output_116_sva_1_mx0, state_output_117_sva_1_mx0, state_output_118_sva_1_mx0,
      state_output_119_sva_1_mx0, state_output_120_sva_1_mx0, state_output_121_sva_1_mx0,
      state_output_122_sva_1_mx0, state_output_123_sva_1_mx0, state_output_124_sva_1_mx0,
      state_output_125_sva_1_mx0, state_output_126_sva_1_mx0, state_output_127_sva_1_mx0,
      operator_ac_int_16_false_1_false_3_acc_nl);
  assign mux_nl = MUX_s_1_2_2(original_rsci_idat, aqed_in_if_issue_dup_aif_1_aif_equal_tmp,
      state_orig_issued_sva);
  assign nl_state_in_count_sva  = state_in_count_sva + 16'b0000000000000001;

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_128_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [15:0] input_56;
    input [15:0] input_57;
    input [15:0] input_58;
    input [15:0] input_59;
    input [15:0] input_60;
    input [15:0] input_61;
    input [15:0] input_62;
    input [15:0] input_63;
    input [15:0] input_64;
    input [15:0] input_65;
    input [15:0] input_66;
    input [15:0] input_67;
    input [15:0] input_68;
    input [15:0] input_69;
    input [15:0] input_70;
    input [15:0] input_71;
    input [15:0] input_72;
    input [15:0] input_73;
    input [15:0] input_74;
    input [15:0] input_75;
    input [15:0] input_76;
    input [15:0] input_77;
    input [15:0] input_78;
    input [15:0] input_79;
    input [15:0] input_80;
    input [15:0] input_81;
    input [15:0] input_82;
    input [15:0] input_83;
    input [15:0] input_84;
    input [15:0] input_85;
    input [15:0] input_86;
    input [15:0] input_87;
    input [15:0] input_88;
    input [15:0] input_89;
    input [15:0] input_90;
    input [15:0] input_91;
    input [15:0] input_92;
    input [15:0] input_93;
    input [15:0] input_94;
    input [15:0] input_95;
    input [15:0] input_96;
    input [15:0] input_97;
    input [15:0] input_98;
    input [15:0] input_99;
    input [15:0] input_100;
    input [15:0] input_101;
    input [15:0] input_102;
    input [15:0] input_103;
    input [15:0] input_104;
    input [15:0] input_105;
    input [15:0] input_106;
    input [15:0] input_107;
    input [15:0] input_108;
    input [15:0] input_109;
    input [15:0] input_110;
    input [15:0] input_111;
    input [15:0] input_112;
    input [15:0] input_113;
    input [15:0] input_114;
    input [15:0] input_115;
    input [15:0] input_116;
    input [15:0] input_117;
    input [15:0] input_118;
    input [15:0] input_119;
    input [15:0] input_120;
    input [15:0] input_121;
    input [15:0] input_122;
    input [15:0] input_123;
    input [15:0] input_124;
    input [15:0] input_125;
    input [15:0] input_126;
    input [15:0] input_127;
    input [6:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      7'b1111101 : begin
        result = input_125;
      end
      7'b1111110 : begin
        result = input_126;
      end
      default : begin
        result = input_127;
      end
    endcase
    MUX_v_16_128_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] conv_u2u_1_7 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_7 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    aqed_top
// ------------------------------------------------------------------


module aqed_top (
  clk, clk_en, reset, bmc_in_rsc_dat, bmc_v_rsc_dat, original_rsc_dat, duplicate_rsc_dat,
      acc_out_rsc_dat, acc_out_v_rsc_dat, acc_out_rdy_rsc_dat, return_aqed_out_rsc_dat,
      return_aqed_out_v_rsc_dat, return_qed_done_rsc_dat, return_qed_check_rsc_dat,
      return_orig_issued_rsc_dat, return_orig_done_rsc_dat
);
  input clk;
  input clk_en;
  input reset;
  input [15:0] bmc_in_rsc_dat;
  input bmc_v_rsc_dat;
  input original_rsc_dat;
  input duplicate_rsc_dat;
  input [15:0] acc_out_rsc_dat;
  input acc_out_v_rsc_dat;
  input acc_out_rdy_rsc_dat;
  output [15:0] return_aqed_out_rsc_dat;
  output return_aqed_out_v_rsc_dat;
  output return_qed_done_rsc_dat;
  output return_qed_check_rsc_dat;
  output return_orig_issued_rsc_dat;
  output return_orig_done_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  aqed_top_core aqed_top_core_inst (
      .clk(clk),
      .clk_en(clk_en),
      .reset(reset),
      .bmc_in_rsc_dat(bmc_in_rsc_dat),
      .bmc_v_rsc_dat(bmc_v_rsc_dat),
      .original_rsc_dat(original_rsc_dat),
      .duplicate_rsc_dat(duplicate_rsc_dat),
      .acc_out_rsc_dat(acc_out_rsc_dat),
      .acc_out_v_rsc_dat(acc_out_v_rsc_dat),
      .acc_out_rdy_rsc_dat(acc_out_rdy_rsc_dat),
      .return_aqed_out_rsc_dat(return_aqed_out_rsc_dat),
      .return_aqed_out_v_rsc_dat(return_aqed_out_v_rsc_dat),
      .return_qed_done_rsc_dat(return_qed_done_rsc_dat),
      .return_qed_check_rsc_dat(return_qed_check_rsc_dat),
      .return_orig_issued_rsc_dat(return_orig_issued_rsc_dat),
      .return_orig_done_rsc_dat(return_orig_done_rsc_dat)
    );
endmodule



